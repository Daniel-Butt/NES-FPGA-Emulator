library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


PACKAGE ROMS IS

	type OAM_REG_ARRAY is array (0 to 255) of std_logic_vector(7 downto 0); -- 64 sprite registers, 4 bytes each
	
   constant OAM_REGS_TEST : OAM_REG_ARRAY := (others=>(others=>'0'));
--	constant OAM_REGS_TEST : OAM_REG_ARRAY := (	x"8C",x"02",x"40",x"37",x"94",x"03",x"40",x"37",x"8C",x"00",x"40",x"3F",x"94",x"01",x"40",x"3F",
--																x"C5",x"9A",x"42",x"8D",x"CD",x"9B",x"42",x"8D",x"C5",x"98",x"42",x"95",x"CD",x"99",x"42",x"95",
--																x"C0",x"9E",x"42",x"5C",x"C8",x"9F",x"42",x"5C",x"C0",x"9C",x"42",x"64",x"C8",x"9D",x"42",x"64",
--																x"4D",x"8C",x"03",x"D5",x"55",x"8D",x"03",x"D5",x"4D",x"8E",x"03",x"DD",x"55",x"8F",x"03",x"DD",
--																x"8B",x"88",x"03",x"9E",x"93",x"89",x"03",x"9E",x"8B",x"8A",x"03",x"A6",x"93",x"8B",x"03",x"A6",
--																x"51",x"88",x"03",x"65",x"59",x"89",x"03",x"65",x"51",x"8A",x"03",x"6D",x"59",x"8B",x"03",x"6D",
--																x"32",x"8C",x"03",x"58",x"3A",x"8D",x"03",x"58",x"32",x"8E",x"03",x"60",x"3A",x"8F",x"03",x"60",
--																x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",
--																x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",
--																x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",
--																x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",
--																x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",x"FF",x"00",x"03",x"00",
--																x"FF",x"D2",x"01",x"BA",x"FF",x"D4",x"01",x"C2",x"FF",x"00",x"01",x"00",x"FF",x"00",x"01",x"00",
--																x"FF",x"F6",x"43",x"98",x"FF",x"F7",x"43",x"98",x"46",x"F6",x"03",x"20",x"4E",x"F7",x"03",x"20",
--																x"C0",x"FC",x"02",x"20",x"C0",x"FD",x"02",x"28",x"18",x"D5",x"01",x"50",x"18",x"D6",x"01",x"58",
--																x"20",x"DB",x"01",x"50",x"28",x"DC",x"01",x"50",x"20",x"DD",x"01",x"58",x"28",x"DE",x"01",x"58");

	type CHR_ROM_ARRAY is array (0 to 8191) of std_logic_vector(7 downto 0);
	
--	constant CHR_ROM_TEST_INIT : CHR_ROM_ARRAY := (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"FF",x"80",x"80",x"00",x"00",x"00",x"80",x"80",x"FF",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
--															x"01",x"01",x"FF",x"01",x"01",x"00",x"00",x"00",x"01",x"01",x"FF",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"FE",x"00",x"C0",x"C0",x"FE",x"7C",x"00",x"7C",x"FE",x"00",x"C0",x"C0",x"FE",x"7C",x"00",x"FE",x"FE",x"00",x"F0",x"C0",x"FE",x"FE",x"00",x"FE",x"FE",x"00",x"F0",x"C0",x"FE",x"FE",x"00",
--															x"C6",x"C6",x"02",x"FE",x"C6",x"C6",x"C6",x"00",x"C6",x"C6",x"02",x"FE",x"C6",x"C6",x"C6",x"00",x"CC",x"D8",x"00",x"F0",x"D8",x"CC",x"C6",x"00",x"CC",x"D8",x"00",x"F0",x"D8",x"CC",x"C6",x"00",x"C6",x"EE",x"02",x"D6",x"C6",x"C6",x"C6",x"00",x"C6",x"EE",x"02",x"D6",x"C6",x"C6",x"C6",x"00",x"C6",x"C6",x"02",x"D6",x"CE",x"C6",x"C6",x"00",x"C6",x"C6",x"02",x"D6",x"CE",x"C6",x"C6",x"00",
--															x"7C",x"FE",x"02",x"C6",x"C6",x"FE",x"7C",x"00",x"7C",x"FE",x"02",x"C6",x"C6",x"FE",x"7C",x"00",x"FC",x"FE",x"02",x"FC",x"C0",x"C0",x"C0",x"00",x"FC",x"FE",x"02",x"FC",x"C0",x"C0",x"C0",x"00",x"CC",x"CC",x"00",x"78",x"30",x"30",x"30",x"00",x"CC",x"CC",x"00",x"78",x"30",x"30",x"30",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",
--															x"FC",x"FE",x"02",x"06",x"1C",x"70",x"FE",x"00",x"FC",x"FE",x"02",x"06",x"1C",x"70",x"FE",x"00",x"FC",x"FE",x"02",x"3C",x"3C",x"02",x"FE",x"00",x"FC",x"FE",x"02",x"3C",x"3C",x"02",x"FE",x"00",x"18",x"18",x"D8",x"D8",x"FE",x"18",x"18",x"00",x"18",x"18",x"D8",x"D8",x"FE",x"18",x"18",x"00",x"FE",x"FE",x"00",x"80",x"FC",x"06",x"FE",x"00",x"FE",x"FE",x"00",x"80",x"FC",x"06",x"FE",x"00",
--															x"7C",x"FE",x"00",x"C0",x"FC",x"C6",x"FE",x"00",x"7C",x"FE",x"00",x"C0",x"FC",x"C6",x"FE",x"00",x"FE",x"FE",x"06",x"0C",x"18",x"10",x"30",x"00",x"FE",x"FE",x"06",x"0C",x"18",x"10",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"33",x"33",x"66",x"00",x"00",x"00",x"00",x"00",x"33",x"33",x"66",x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"FF",x"66",x"FF",x"66",x"66",x"00",x"66",x"66",x"FF",x"66",x"FF",x"66",x"66",x"00",
--															x"18",x"3E",x"60",x"3C",x"06",x"7C",x"18",x"00",x"18",x"3E",x"60",x"3C",x"06",x"7C",x"18",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"46",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"46",x"00",x"3C",x"66",x"3C",x"38",x"67",x"66",x"3F",x"00",x"3C",x"66",x"3C",x"38",x"67",x"66",x"3F",x"00",x"0C",x"0C",x"18",x"00",x"00",x"00",x"00",x"00",x"0C",x"0C",x"18",x"00",x"00",x"00",x"00",x"00",
--															x"0C",x"18",x"30",x"30",x"30",x"18",x"0C",x"00",x"0C",x"18",x"30",x"30",x"30",x"18",x"0C",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"18",x"30",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"18",x"30",x"00",x"00",x"66",x"3C",x"FF",x"3C",x"66",x"00",x"00",x"00",x"66",x"3C",x"FF",x"3C",x"66",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"6E",x"3B",x"00",x"00",x"00",x"00",x"00",x"00",x"6E",x"3B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"03",x"06",x"0C",x"18",x"30",x"60",x"00",x"00",x"03",x"06",x"0C",x"18",x"30",x"60",x"00",
--															x"3E",x"63",x"67",x"6B",x"73",x"63",x"3E",x"00",x"3E",x"63",x"67",x"6B",x"73",x"63",x"3E",x"00",x"0C",x"1C",x"0C",x"0C",x"0C",x"0C",x"3F",x"00",x"0C",x"1C",x"0C",x"0C",x"0C",x"0C",x"3F",x"00",x"3E",x"63",x"63",x"0E",x"38",x"63",x"7F",x"00",x"3E",x"63",x"63",x"0E",x"38",x"63",x"7F",x"00",x"3E",x"63",x"63",x"0E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"63",x"0E",x"63",x"63",x"3E",x"00",
--															x"06",x"0E",x"1E",x"26",x"7F",x"06",x"06",x"00",x"06",x"0E",x"1E",x"26",x"7F",x"06",x"06",x"00",x"7F",x"63",x"60",x"7E",x"03",x"63",x"3E",x"00",x"7F",x"63",x"60",x"7E",x"03",x"63",x"3E",x"00",x"3E",x"63",x"60",x"7E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"60",x"7E",x"63",x"63",x"3E",x"00",x"7F",x"63",x"06",x"0C",x"18",x"18",x"3C",x"00",x"7F",x"63",x"06",x"0C",x"18",x"18",x"3C",x"00",
--															x"3E",x"63",x"63",x"3E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"63",x"3E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"63",x"3F",x"03",x"63",x"3E",x"00",x"3E",x"63",x"63",x"3F",x"03",x"63",x"3E",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"30",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"30",
--															x"0E",x"18",x"30",x"60",x"30",x"18",x"0E",x"00",x"0E",x"18",x"30",x"60",x"30",x"18",x"0E",x"00",x"00",x"00",x"7E",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"7E",x"00",x"00",x"00",x"70",x"18",x"0C",x"06",x"0C",x"18",x"70",x"00",x"70",x"18",x"0C",x"06",x"0C",x"18",x"70",x"00",x"7E",x"63",x"03",x"06",x"1C",x"00",x"18",x"18",x"7E",x"63",x"03",x"06",x"1C",x"00",x"18",x"18",
--															x"7C",x"C6",x"CE",x"EE",x"E0",x"E6",x"7C",x"00",x"7C",x"C6",x"CE",x"EE",x"E0",x"E6",x"7C",x"00",x"1C",x"36",x"63",x"7F",x"63",x"63",x"63",x"00",x"1C",x"36",x"63",x"7F",x"63",x"63",x"63",x"00",x"6E",x"73",x"63",x"7E",x"63",x"63",x"7E",x"00",x"6E",x"73",x"63",x"7E",x"63",x"63",x"7E",x"00",x"1E",x"33",x"60",x"60",x"60",x"33",x"1E",x"00",x"1E",x"33",x"60",x"60",x"60",x"33",x"1E",x"00",
--															x"6C",x"76",x"63",x"63",x"63",x"66",x"7C",x"00",x"6C",x"76",x"63",x"63",x"63",x"66",x"7C",x"00",x"7F",x"31",x"30",x"3C",x"30",x"31",x"7F",x"00",x"7F",x"31",x"30",x"3C",x"30",x"31",x"7F",x"00",x"7F",x"31",x"30",x"3C",x"30",x"30",x"78",x"00",x"7F",x"31",x"30",x"3C",x"30",x"30",x"78",x"00",x"1E",x"33",x"60",x"67",x"63",x"37",x"1D",x"00",x"1E",x"33",x"60",x"67",x"63",x"37",x"1D",x"00",
--															x"63",x"63",x"63",x"7F",x"63",x"63",x"63",x"00",x"63",x"63",x"63",x"7F",x"63",x"63",x"63",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"1F",x"06",x"06",x"06",x"06",x"66",x"3C",x"00",x"1F",x"06",x"06",x"06",x"06",x"66",x"3C",x"00",x"66",x"66",x"6C",x"78",x"6C",x"67",x"63",x"00",x"66",x"66",x"6C",x"78",x"6C",x"67",x"63",x"00",
--															x"78",x"30",x"60",x"60",x"63",x"63",x"7E",x"00",x"78",x"30",x"60",x"60",x"63",x"63",x"7E",x"00",x"63",x"77",x"7F",x"6B",x"63",x"63",x"63",x"00",x"63",x"77",x"7F",x"6B",x"63",x"63",x"63",x"00",x"63",x"73",x"7B",x"6F",x"67",x"63",x"63",x"00",x"63",x"73",x"7B",x"6F",x"67",x"63",x"63",x"00",x"1C",x"36",x"63",x"63",x"63",x"36",x"1C",x"00",x"1C",x"36",x"63",x"63",x"63",x"36",x"1C",x"00",
--															x"6E",x"73",x"63",x"7E",x"60",x"60",x"60",x"00",x"6E",x"73",x"63",x"7E",x"60",x"60",x"60",x"00",x"1C",x"36",x"63",x"6B",x"67",x"36",x"1D",x"00",x"1C",x"36",x"63",x"6B",x"67",x"36",x"1D",x"00",x"6E",x"73",x"63",x"7E",x"6C",x"67",x"63",x"00",x"6E",x"73",x"63",x"7E",x"6C",x"67",x"63",x"00",x"3E",x"63",x"60",x"3E",x"03",x"63",x"3E",x"00",x"3E",x"63",x"60",x"3E",x"03",x"63",x"3E",x"00",
--															x"7E",x"5A",x"18",x"18",x"18",x"18",x"3C",x"00",x"7E",x"5A",x"18",x"18",x"18",x"18",x"3C",x"00",x"73",x"33",x"63",x"63",x"63",x"76",x"3C",x"00",x"73",x"33",x"63",x"63",x"63",x"76",x"3C",x"00",x"73",x"33",x"63",x"63",x"66",x"3C",x"18",x"00",x"73",x"33",x"63",x"63",x"66",x"3C",x"18",x"00",x"73",x"33",x"63",x"6B",x"7F",x"77",x"63",x"00",x"73",x"33",x"63",x"6B",x"7F",x"77",x"63",x"00",
--															x"63",x"63",x"36",x"1C",x"36",x"63",x"63",x"00",x"63",x"63",x"36",x"1C",x"36",x"63",x"63",x"00",x"33",x"63",x"63",x"36",x"1C",x"78",x"70",x"00",x"33",x"63",x"63",x"36",x"1C",x"78",x"70",x"00",x"7F",x"63",x"06",x"1C",x"33",x"63",x"7E",x"00",x"7F",x"63",x"06",x"1C",x"33",x"63",x"7E",x"00",x"3C",x"30",x"30",x"30",x"30",x"30",x"3C",x"00",x"3C",x"30",x"30",x"30",x"30",x"30",x"3C",x"00",
--															x"40",x"60",x"30",x"18",x"0C",x"06",x"02",x"00",x"40",x"60",x"30",x"18",x"0C",x"06",x"02",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
--															x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"63",x"63",x"67",x"3B",x"00",x"00",x"00",x"3F",x"63",x"63",x"67",x"3B",x"00",x"60",x"60",x"6E",x"73",x"63",x"63",x"3E",x"00",x"60",x"60",x"6E",x"73",x"63",x"63",x"3E",x"00",x"00",x"00",x"3E",x"63",x"60",x"63",x"3E",x"00",x"00",x"00",x"3E",x"63",x"60",x"63",x"3E",x"00",
--															x"03",x"03",x"3B",x"67",x"63",x"63",x"3E",x"00",x"03",x"03",x"3B",x"67",x"63",x"63",x"3E",x"00",x"00",x"00",x"3E",x"61",x"7F",x"60",x"3E",x"00",x"00",x"00",x"3E",x"61",x"7F",x"60",x"3E",x"00",x"0E",x"18",x"18",x"3C",x"18",x"18",x"3C",x"00",x"0E",x"18",x"18",x"3C",x"18",x"18",x"3C",x"00",x"00",x"00",x"3E",x"60",x"63",x"63",x"3D",x"00",x"00",x"00",x"3E",x"60",x"63",x"63",x"3D",x"00",
--															x"60",x"60",x"6E",x"73",x"63",x"66",x"67",x"00",x"60",x"60",x"6E",x"73",x"63",x"66",x"67",x"00",x"00",x"00",x"1E",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"1E",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"3F",x"06",x"06",x"06",x"66",x"3C",x"00",x"00",x"3F",x"06",x"06",x"06",x"66",x"3C",x"60",x"60",x"66",x"6E",x"7C",x"67",x"63",x"00",x"60",x"60",x"66",x"6E",x"7C",x"67",x"63",x"00",
--															x"1C",x"0C",x"0C",x"0C",x"0C",x"0C",x"1E",x"00",x"1C",x"0C",x"0C",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"6E",x"7F",x"6B",x"62",x"67",x"00",x"00",x"00",x"6E",x"7F",x"6B",x"62",x"67",x"00",x"00",x"00",x"6E",x"73",x"63",x"66",x"67",x"00",x"00",x"00",x"6E",x"73",x"63",x"66",x"67",x"00",x"00",x"00",x"3E",x"63",x"63",x"63",x"3E",x"00",x"00",x"00",x"3E",x"63",x"63",x"63",x"3E",x"00",
--															x"00",x"00",x"3E",x"63",x"73",x"6E",x"60",x"60",x"00",x"00",x"3E",x"63",x"73",x"6E",x"60",x"60",x"00",x"00",x"3E",x"63",x"67",x"3B",x"03",x"03",x"00",x"00",x"3E",x"63",x"67",x"3B",x"03",x"03",x"00",x"00",x"6E",x"73",x"63",x"7E",x"63",x"00",x"00",x"00",x"6E",x"73",x"63",x"7E",x"63",x"00",x"00",x"00",x"3E",x"71",x"1C",x"47",x"3E",x"00",x"00",x"00",x"3E",x"71",x"1C",x"47",x"3E",x"00",
--															x"06",x"0C",x"3F",x"18",x"18",x"1B",x"0E",x"00",x"06",x"0C",x"3F",x"18",x"18",x"1B",x"0E",x"00",x"00",x"00",x"73",x"33",x"63",x"67",x"3B",x"00",x"00",x"00",x"73",x"33",x"63",x"67",x"3B",x"00",x"00",x"00",x"73",x"33",x"63",x"66",x"3C",x"00",x"00",x"00",x"73",x"33",x"63",x"66",x"3C",x"00",x"00",x"00",x"63",x"6B",x"7F",x"77",x"63",x"00",x"00",x"00",x"63",x"6B",x"7F",x"77",x"63",x"00",
--															x"00",x"00",x"63",x"36",x"1C",x"36",x"63",x"00",x"00",x"00",x"63",x"36",x"1C",x"36",x"63",x"00",x"00",x"00",x"33",x"63",x"63",x"3F",x"03",x"3E",x"00",x"00",x"33",x"63",x"63",x"3F",x"03",x"3E",x"00",x"00",x"7F",x"0E",x"1C",x"38",x"7F",x"00",x"00",x"00",x"7F",x"0E",x"1C",x"38",x"7F",x"00",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
--	
	
	
	constant NES_TEST_CHR_ROM : CHR_ROM_ARRAY := (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"FF",x"80",x"80",x"00",x"00",x"00",x"80",x"80",x"FF",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
																	x"01",x"01",x"FF",x"01",x"01",x"00",x"00",x"00",x"01",x"01",x"FF",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"FE",x"00",x"C0",x"C0",x"FE",x"7C",x"00",x"7C",x"FE",x"00",x"C0",x"C0",x"FE",x"7C",x"00",x"FE",x"FE",x"00",x"F0",x"C0",x"FE",x"FE",x"00",x"FE",x"FE",x"00",x"F0",x"C0",x"FE",x"FE",x"00",
																	x"C6",x"C6",x"02",x"FE",x"C6",x"C6",x"C6",x"00",x"C6",x"C6",x"02",x"FE",x"C6",x"C6",x"C6",x"00",x"CC",x"D8",x"00",x"F0",x"D8",x"CC",x"C6",x"00",x"CC",x"D8",x"00",x"F0",x"D8",x"CC",x"C6",x"00",x"C6",x"EE",x"02",x"D6",x"C6",x"C6",x"C6",x"00",x"C6",x"EE",x"02",x"D6",x"C6",x"C6",x"C6",x"00",x"C6",x"C6",x"02",x"D6",x"CE",x"C6",x"C6",x"00",x"C6",x"C6",x"02",x"D6",x"CE",x"C6",x"C6",x"00",
																	x"7C",x"FE",x"02",x"C6",x"C6",x"FE",x"7C",x"00",x"7C",x"FE",x"02",x"C6",x"C6",x"FE",x"7C",x"00",x"FC",x"FE",x"02",x"FC",x"C0",x"C0",x"C0",x"00",x"FC",x"FE",x"02",x"FC",x"C0",x"C0",x"C0",x"00",x"CC",x"CC",x"00",x"78",x"30",x"30",x"30",x"00",x"CC",x"CC",x"00",x"78",x"30",x"30",x"30",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",
																	x"FC",x"FE",x"02",x"06",x"1C",x"70",x"FE",x"00",x"FC",x"FE",x"02",x"06",x"1C",x"70",x"FE",x"00",x"FC",x"FE",x"02",x"3C",x"3C",x"02",x"FE",x"00",x"FC",x"FE",x"02",x"3C",x"3C",x"02",x"FE",x"00",x"18",x"18",x"D8",x"D8",x"FE",x"18",x"18",x"00",x"18",x"18",x"D8",x"D8",x"FE",x"18",x"18",x"00",x"FE",x"FE",x"00",x"80",x"FC",x"06",x"FE",x"00",x"FE",x"FE",x"00",x"80",x"FC",x"06",x"FE",x"00",
																	x"7C",x"FE",x"00",x"C0",x"FC",x"C6",x"FE",x"00",x"7C",x"FE",x"00",x"C0",x"FC",x"C6",x"FE",x"00",x"FE",x"FE",x"06",x"0C",x"18",x"10",x"30",x"00",x"FE",x"FE",x"06",x"0C",x"18",x"10",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"33",x"33",x"66",x"00",x"00",x"00",x"00",x"00",x"33",x"33",x"66",x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"FF",x"66",x"FF",x"66",x"66",x"00",x"66",x"66",x"FF",x"66",x"FF",x"66",x"66",x"00",
																	x"18",x"3E",x"60",x"3C",x"06",x"7C",x"18",x"00",x"18",x"3E",x"60",x"3C",x"06",x"7C",x"18",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"46",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"46",x"00",x"3C",x"66",x"3C",x"38",x"67",x"66",x"3F",x"00",x"3C",x"66",x"3C",x"38",x"67",x"66",x"3F",x"00",x"0C",x"0C",x"18",x"00",x"00",x"00",x"00",x"00",x"0C",x"0C",x"18",x"00",x"00",x"00",x"00",x"00",
																	x"0C",x"18",x"30",x"30",x"30",x"18",x"0C",x"00",x"0C",x"18",x"30",x"30",x"30",x"18",x"0C",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"18",x"30",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"18",x"30",x"00",x"00",x"66",x"3C",x"FF",x"3C",x"66",x"00",x"00",x"00",x"66",x"3C",x"FF",x"3C",x"66",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"6E",x"3B",x"00",x"00",x"00",x"00",x"00",x"00",x"6E",x"3B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"03",x"06",x"0C",x"18",x"30",x"60",x"00",x"00",x"03",x"06",x"0C",x"18",x"30",x"60",x"00",
																	x"3E",x"63",x"67",x"6B",x"73",x"63",x"3E",x"00",x"3E",x"63",x"67",x"6B",x"73",x"63",x"3E",x"00",x"0C",x"1C",x"0C",x"0C",x"0C",x"0C",x"3F",x"00",x"0C",x"1C",x"0C",x"0C",x"0C",x"0C",x"3F",x"00",x"3E",x"63",x"63",x"0E",x"38",x"63",x"7F",x"00",x"3E",x"63",x"63",x"0E",x"38",x"63",x"7F",x"00",x"3E",x"63",x"63",x"0E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"63",x"0E",x"63",x"63",x"3E",x"00",
																	x"06",x"0E",x"1E",x"26",x"7F",x"06",x"06",x"00",x"06",x"0E",x"1E",x"26",x"7F",x"06",x"06",x"00",x"7F",x"63",x"60",x"7E",x"03",x"63",x"3E",x"00",x"7F",x"63",x"60",x"7E",x"03",x"63",x"3E",x"00",x"3E",x"63",x"60",x"7E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"60",x"7E",x"63",x"63",x"3E",x"00",x"7F",x"63",x"06",x"0C",x"18",x"18",x"3C",x"00",x"7F",x"63",x"06",x"0C",x"18",x"18",x"3C",x"00",
																	x"3E",x"63",x"63",x"3E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"63",x"3E",x"63",x"63",x"3E",x"00",x"3E",x"63",x"63",x"3F",x"03",x"63",x"3E",x"00",x"3E",x"63",x"63",x"3F",x"03",x"63",x"3E",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"30",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"30",
																	x"0E",x"18",x"30",x"60",x"30",x"18",x"0E",x"00",x"0E",x"18",x"30",x"60",x"30",x"18",x"0E",x"00",x"00",x"00",x"7E",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"7E",x"00",x"00",x"00",x"70",x"18",x"0C",x"06",x"0C",x"18",x"70",x"00",x"70",x"18",x"0C",x"06",x"0C",x"18",x"70",x"00",x"7E",x"63",x"03",x"06",x"1C",x"00",x"18",x"18",x"7E",x"63",x"03",x"06",x"1C",x"00",x"18",x"18",
																	x"7C",x"C6",x"CE",x"EE",x"E0",x"E6",x"7C",x"00",x"7C",x"C6",x"CE",x"EE",x"E0",x"E6",x"7C",x"00",x"1C",x"36",x"63",x"7F",x"63",x"63",x"63",x"00",x"1C",x"36",x"63",x"7F",x"63",x"63",x"63",x"00",x"6E",x"73",x"63",x"7E",x"63",x"63",x"7E",x"00",x"6E",x"73",x"63",x"7E",x"63",x"63",x"7E",x"00",x"1E",x"33",x"60",x"60",x"60",x"33",x"1E",x"00",x"1E",x"33",x"60",x"60",x"60",x"33",x"1E",x"00",
																	x"6C",x"76",x"63",x"63",x"63",x"66",x"7C",x"00",x"6C",x"76",x"63",x"63",x"63",x"66",x"7C",x"00",x"7F",x"31",x"30",x"3C",x"30",x"31",x"7F",x"00",x"7F",x"31",x"30",x"3C",x"30",x"31",x"7F",x"00",x"7F",x"31",x"30",x"3C",x"30",x"30",x"78",x"00",x"7F",x"31",x"30",x"3C",x"30",x"30",x"78",x"00",x"1E",x"33",x"60",x"67",x"63",x"37",x"1D",x"00",x"1E",x"33",x"60",x"67",x"63",x"37",x"1D",x"00",
																	x"63",x"63",x"63",x"7F",x"63",x"63",x"63",x"00",x"63",x"63",x"63",x"7F",x"63",x"63",x"63",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"1F",x"06",x"06",x"06",x"06",x"66",x"3C",x"00",x"1F",x"06",x"06",x"06",x"06",x"66",x"3C",x"00",x"66",x"66",x"6C",x"78",x"6C",x"67",x"63",x"00",x"66",x"66",x"6C",x"78",x"6C",x"67",x"63",x"00",
																	x"78",x"30",x"60",x"60",x"63",x"63",x"7E",x"00",x"78",x"30",x"60",x"60",x"63",x"63",x"7E",x"00",x"63",x"77",x"7F",x"6B",x"63",x"63",x"63",x"00",x"63",x"77",x"7F",x"6B",x"63",x"63",x"63",x"00",x"63",x"73",x"7B",x"6F",x"67",x"63",x"63",x"00",x"63",x"73",x"7B",x"6F",x"67",x"63",x"63",x"00",x"1C",x"36",x"63",x"63",x"63",x"36",x"1C",x"00",x"1C",x"36",x"63",x"63",x"63",x"36",x"1C",x"00",
																	x"6E",x"73",x"63",x"7E",x"60",x"60",x"60",x"00",x"6E",x"73",x"63",x"7E",x"60",x"60",x"60",x"00",x"1C",x"36",x"63",x"6B",x"67",x"36",x"1D",x"00",x"1C",x"36",x"63",x"6B",x"67",x"36",x"1D",x"00",x"6E",x"73",x"63",x"7E",x"6C",x"67",x"63",x"00",x"6E",x"73",x"63",x"7E",x"6C",x"67",x"63",x"00",x"3E",x"63",x"60",x"3E",x"03",x"63",x"3E",x"00",x"3E",x"63",x"60",x"3E",x"03",x"63",x"3E",x"00",
																	x"7E",x"5A",x"18",x"18",x"18",x"18",x"3C",x"00",x"7E",x"5A",x"18",x"18",x"18",x"18",x"3C",x"00",x"73",x"33",x"63",x"63",x"63",x"76",x"3C",x"00",x"73",x"33",x"63",x"63",x"63",x"76",x"3C",x"00",x"73",x"33",x"63",x"63",x"66",x"3C",x"18",x"00",x"73",x"33",x"63",x"63",x"66",x"3C",x"18",x"00",x"73",x"33",x"63",x"6B",x"7F",x"77",x"63",x"00",x"73",x"33",x"63",x"6B",x"7F",x"77",x"63",x"00",
																	x"63",x"63",x"36",x"1C",x"36",x"63",x"63",x"00",x"63",x"63",x"36",x"1C",x"36",x"63",x"63",x"00",x"33",x"63",x"63",x"36",x"1C",x"78",x"70",x"00",x"33",x"63",x"63",x"36",x"1C",x"78",x"70",x"00",x"7F",x"63",x"06",x"1C",x"33",x"63",x"7E",x"00",x"7F",x"63",x"06",x"1C",x"33",x"63",x"7E",x"00",x"3C",x"30",x"30",x"30",x"30",x"30",x"3C",x"00",x"3C",x"30",x"30",x"30",x"30",x"30",x"3C",x"00",
																	x"40",x"60",x"30",x"18",x"0C",x"06",x"02",x"00",x"40",x"60",x"30",x"18",x"0C",x"06",x"02",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
																	x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"63",x"63",x"67",x"3B",x"00",x"00",x"00",x"3F",x"63",x"63",x"67",x"3B",x"00",x"60",x"60",x"6E",x"73",x"63",x"63",x"3E",x"00",x"60",x"60",x"6E",x"73",x"63",x"63",x"3E",x"00",x"00",x"00",x"3E",x"63",x"60",x"63",x"3E",x"00",x"00",x"00",x"3E",x"63",x"60",x"63",x"3E",x"00",
																	x"03",x"03",x"3B",x"67",x"63",x"63",x"3E",x"00",x"03",x"03",x"3B",x"67",x"63",x"63",x"3E",x"00",x"00",x"00",x"3E",x"61",x"7F",x"60",x"3E",x"00",x"00",x"00",x"3E",x"61",x"7F",x"60",x"3E",x"00",x"0E",x"18",x"18",x"3C",x"18",x"18",x"3C",x"00",x"0E",x"18",x"18",x"3C",x"18",x"18",x"3C",x"00",x"00",x"00",x"3E",x"60",x"63",x"63",x"3D",x"00",x"00",x"00",x"3E",x"60",x"63",x"63",x"3D",x"00",
																	x"60",x"60",x"6E",x"73",x"63",x"66",x"67",x"00",x"60",x"60",x"6E",x"73",x"63",x"66",x"67",x"00",x"00",x"00",x"1E",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"1E",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"3F",x"06",x"06",x"06",x"66",x"3C",x"00",x"00",x"3F",x"06",x"06",x"06",x"66",x"3C",x"60",x"60",x"66",x"6E",x"7C",x"67",x"63",x"00",x"60",x"60",x"66",x"6E",x"7C",x"67",x"63",x"00",
																	x"1C",x"0C",x"0C",x"0C",x"0C",x"0C",x"1E",x"00",x"1C",x"0C",x"0C",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",x"6E",x"7F",x"6B",x"62",x"67",x"00",x"00",x"00",x"6E",x"7F",x"6B",x"62",x"67",x"00",x"00",x"00",x"6E",x"73",x"63",x"66",x"67",x"00",x"00",x"00",x"6E",x"73",x"63",x"66",x"67",x"00",x"00",x"00",x"3E",x"63",x"63",x"63",x"3E",x"00",x"00",x"00",x"3E",x"63",x"63",x"63",x"3E",x"00",
																	x"00",x"00",x"3E",x"63",x"73",x"6E",x"60",x"60",x"00",x"00",x"3E",x"63",x"73",x"6E",x"60",x"60",x"00",x"00",x"3E",x"63",x"67",x"3B",x"03",x"03",x"00",x"00",x"3E",x"63",x"67",x"3B",x"03",x"03",x"00",x"00",x"6E",x"73",x"63",x"7E",x"63",x"00",x"00",x"00",x"6E",x"73",x"63",x"7E",x"63",x"00",x"00",x"00",x"3E",x"71",x"1C",x"47",x"3E",x"00",x"00",x"00",x"3E",x"71",x"1C",x"47",x"3E",x"00",
																	x"06",x"0C",x"3F",x"18",x"18",x"1B",x"0E",x"00",x"06",x"0C",x"3F",x"18",x"18",x"1B",x"0E",x"00",x"00",x"00",x"73",x"33",x"63",x"67",x"3B",x"00",x"00",x"00",x"73",x"33",x"63",x"67",x"3B",x"00",x"00",x"00",x"73",x"33",x"63",x"66",x"3C",x"00",x"00",x"00",x"73",x"33",x"63",x"66",x"3C",x"00",x"00",x"00",x"63",x"6B",x"7F",x"77",x"63",x"00",x"00",x"00",x"63",x"6B",x"7F",x"77",x"63",x"00",
																	x"00",x"00",x"63",x"36",x"1C",x"36",x"63",x"00",x"00",x"00",x"63",x"36",x"1C",x"36",x"63",x"00",x"00",x"00",x"33",x"63",x"63",x"3F",x"03",x"3E",x"00",x"00",x"33",x"63",x"63",x"3F",x"03",x"3E",x"00",x"00",x"7F",x"0E",x"1C",x"38",x"7F",x"00",x"00",x"00",x"7F",x"0E",x"1C",x"38",x"7F",x"00",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
	
	
	constant FOOTBALL_CHR_ROM : CHR_ROM_ARRAY := (x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00", x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00", x"0C", x"1C", x"0C", x"0C", x"0C", x"0C", x"3F", x"00", x"0C", x"1C", x"0C", x"0C", x"0C", x"0C", x"3F", x"00", x"3E", x"63", x"07", x"1E", x"3C", x"70", x"7F", x"00", x"3E", x"63", x"07", x"1E", x"3C", x"70", x"7F", x"00", x"3F", x"06", x"0C", x"1E", x"03", x"63", x"3E", x"00", x"3F", x"06", x"0C", x"1E", x"03", x"63", x"3E", x"00", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"7E", x"60", x"7E", x"03", x"03", x"63", x"3E", x"00", x"7E", x"60", x"7E", x"03", x"03", x"63", x"3E", x"00", x"1E", x"30", x"60", x"7E", x"63", x"63", x"3E", x"00", x"1E", x"30", x"60", x"7E", x"63", x"63", x"3E", x"00", x"7F", x"63", x"06", x"0C", x"18", x"18", x"18", x"00", x"7F", x"63", x"06", x"0C", x"18", x"18", x"18", x"00", 
															x"3C", x"62", x"72", x"3C", x"4F", x"43", x"3E", x"00", x"3C", x"62", x"72", x"3C", x"4F", x"43", x"3E", x"00", x"3E", x"63", x"63", x"3F", x"03", x"06", x"3C", x"00", x"3E", x"63", x"63", x"3F", x"03", x"06", x"3C", x"00", x"1C", x"36", x"63", x"63", x"7F", x"63", x"63", x"00", x"1C", x"36", x"63", x"63", x"7F", x"63", x"63", x"00", x"7E", x"63", x"63", x"7E", x"63", x"63", x"7E", x"00", x"7E", x"63", x"63", x"7E", x"63", x"63", x"7E", x"00", x"1E", x"33", x"60", x"60", x"60", x"33", x"1E", x"00", x"1E", x"33", x"60", x"60", x"60", x"33", x"1E", x"00", x"7C", x"66", x"63", x"63", x"63", x"66", x"7C", x"00", x"7C", x"66", x"63", x"63", x"63", x"66", x"7C", x"00", x"3F", x"30", x"30", x"3E", x"30", x"30", x"3F", x"00", x"3F", x"30", x"30", x"3E", x"30", x"30", x"3F", x"00", x"7F", x"60", x"60", x"7E", x"60", x"60", x"60", x"00", x"7F", x"60", x"60", x"7E", x"60", x"60", x"60", x"00", 
															x"1F", x"30", x"60", x"67", x"63", x"33", x"1F", x"00", x"1F", x"30", x"60", x"67", x"63", x"33", x"1F", x"00", x"63", x"63", x"63", x"7F", x"63", x"63", x"63", x"00", x"63", x"63", x"63", x"7F", x"63", x"63", x"63", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00", x"03", x"03", x"03", x"03", x"03", x"63", x"3E", x"00", x"03", x"03", x"03", x"03", x"03", x"63", x"3E", x"00", x"63", x"66", x"6C", x"78", x"7C", x"6E", x"67", x"00", x"63", x"66", x"6C", x"78", x"7C", x"6E", x"67", x"00", x"30", x"30", x"30", x"30", x"30", x"30", x"3F", x"00", x"30", x"30", x"30", x"30", x"30", x"30", x"3F", x"00", x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00", x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00", x"63", x"73", x"7B", x"7F", x"6F", x"67", x"63", x"00", x"63", x"73", x"7B", x"7F", x"6F", x"67", x"63", x"00", 
															x"3E", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"3E", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"7E", x"63", x"63", x"63", x"7E", x"60", x"60", x"00", x"7E", x"63", x"63", x"63", x"7E", x"60", x"60", x"00", x"3E", x"63", x"63", x"63", x"6F", x"66", x"3D", x"00", x"3E", x"63", x"63", x"63", x"6F", x"66", x"3D", x"00", x"7E", x"63", x"63", x"67", x"7C", x"6E", x"67", x"00", x"7E", x"63", x"63", x"67", x"7C", x"6E", x"67", x"00", x"3C", x"66", x"60", x"3E", x"03", x"63", x"3E", x"00", x"3C", x"66", x"60", x"3E", x"03", x"63", x"3E", x"00", x"3F", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"3F", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"63", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"63", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"63", x"63", x"63", x"77", x"3E", x"1C", x"08", x"00", x"63", x"63", x"63", x"77", x"3E", x"1C", x"08", x"00", 
															x"63", x"63", x"6B", x"7F", x"7F", x"36", x"22", x"00", x"63", x"63", x"6B", x"7F", x"7F", x"36", x"22", x"00", x"63", x"77", x"3E", x"1C", x"3E", x"77", x"63", x"00", x"63", x"77", x"3E", x"1C", x"3E", x"77", x"63", x"00", x"33", x"33", x"12", x"1E", x"0C", x"0C", x"0C", x"00", x"33", x"33", x"12", x"1E", x"0C", x"0C", x"0C", x"00", x"7F", x"07", x"0E", x"1C", x"38", x"70", x"7F", x"00", x"7F", x"07", x"0E", x"1C", x"38", x"70", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"04", x"04", x"04", x"6F", x"84", x"64", x"14", x"E3", x"04", x"04", x"04", x"6F", x"84", x"64", x"14", x"E3", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"44", x"4A", x"52", x"53", x"4D", x"00", x"40", x"40", x"44", x"4A", x"52", x"53", x"4D", 
															x"00", x"00", x"00", x"64", x"8E", x"64", x"15", x"E2", x"00", x"00", x"00", x"64", x"8E", x"64", x"15", x"E2", x"00", x"82", x"45", x"29", x"2A", x"12", x"13", x"12", x"00", x"82", x"45", x"29", x"2A", x"12", x"13", x"12", x"00", x"8F", x"48", x"48", x"2F", x"29", x"E8", x"28", x"00", x"8F", x"48", x"48", x"2F", x"29", x"E8", x"28", x"00", x"38", x"A4", x"A2", x"22", x"22", x"A4", x"78", x"00", x"38", x"A4", x"A2", x"22", x"22", x"A4", x"78", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"6C", x"5E", x"5C", x"60", x"30", x"01", x"00", x"00", x"0C", x"1E", x"18", x"1C", x"0E", x"3E", x"3E", x"3C", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"76", x"67", x"67", x"06", x"06", x"00", x"00", x"3C", x"76", x"67", x"67", x"60", x"00", x"06", x"07", x"00", x"00", x"18", x"3C", x"00", x"80", x"C2", x"40", x"00", x"00", x"18", x"3C", x"7E", x"7F", x"3C", x"3C", x"3C", x"7E", x"77", x"67", x"66", x"06", x"00", x"00", x"3C", x"7E", x"77", x"07", x"04", x"60", x"06", x"07", x"00", x"18", x"3C", x"04", x"00", x"08", x"0C", x"07", x"00", x"18", x"3C", x"7C", x"7C", x"F4", x"F0", x"F8", x"3C", x"7E", x"66", x"66", x"C4", x"80", x"00", x"00", x"3C", x"7E", x"66", x"60", x"00", x"06", x"C0", x"00", x"7C", x"3C", x"3C", x"6C", x"4C", x"08", x"00", x"00", x"7C", x"3C", x"3C", x"0C", x"80", x"40", x"0C", x"00", x"18", x"7C", x"3C", x"00", x"00", x"81", x"81", x"C3", x"18", x"7C", x"1C", x"7E", x"FF", x"7E", x"3C", x"3C", 
															x"3C", x"6C", x"6C", x"CC", x"C6", x"66", x"22", x"00", x"3C", x"6C", x"6C", x"CC", x"C2", x"00", x"00", x"66", x"18", x"3C", x"38", x"18", x"00", x"40", x"C6", x"0C", x"18", x"3C", x"20", x"26", x"7F", x"3F", x"38", x"12", x"3E", x"7E", x"6C", x"D8", x"CC", x"4C", x"04", x"00", x"3E", x"7E", x"6C", x"58", x"04", x"00", x"C2", x"0C", x"0C", x"1E", x"0E", x"00", x"00", x"80", x"E1", x"00", x"0C", x"1E", x"02", x"1E", x"3F", x"3F", x"1E", x"1E", x"3E", x"3C", x"78", x"D8", x"CC", x"66", x"62", x"00", x"3E", x"3C", x"78", x"D8", x"C8", x"00", x"01", x"E6", x"18", x"3C", x"38", x"18", x"00", x"81", x"C3", x"66", x"18", x"3C", x"20", x"66", x"FF", x"7E", x"3C", x"18", x"3E", x"3E", x"6C", x"6C", x"6C", x"66", x"62", x"00", x"3E", x"3E", x"6C", x"6C", x"2C", x"00", x"01", x"E6", x"18", x"3C", x"38", x"18", x"00", x"81", x"81", x"C3", x"18", x"3C", x"20", x"66", x"FF", x"7E", x"7E", x"3C", 
															x"3C", x"3C", x"6C", x"6C", x"6C", x"64", x"24", x"00", x"3C", x"3C", x"6C", x"6C", x"28", x"02", x"02", x"64", x"80", x"C0", x"B0", x"F8", x"80", x"00", x"01", x"00", x"00", x"00", x"30", x"78", x"7E", x"7F", x"3E", x"1E", x"1E", x"3C", x"78", x"38", x"18", x"0C", x"04", x"00", x"1E", x"3C", x"78", x"38", x"78", x"00", x"00", x"0C", x"1E", x"3C", x"3C", x"36", x"32", x"10", x"00", x"00", x"1E", x"3C", x"3C", x"30", x"01", x"02", x"30", x"00", x"3C", x"7E", x"66", x"66", x"43", x"01", x"00", x"00", x"3C", x"7E", x"66", x"26", x"20", x"C0", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0D", x"1F", x"1F", x"0C", x"00", x"80", x"C0", x"40", x"0C", x"1E", x"12", x"33", x"7F", x"7E", x"3E", x"3E", x"0D", x"1F", x"1D", x"0C", x"00", x"80", x"C0", x"60", x"0C", x"1E", x"10", x"33", x"7F", x"7E", x"3E", x"1E", 
															x"0D", x"1F", x"1D", x"0C", x"00", x"C0", x"60", x"30", x"0C", x"1E", x"10", x"33", x"7F", x"3E", x"1E", x"0E", x"0C", x"1E", x"1C", x"0C", x"00", x"81", x"C3", x"46", x"0C", x"1E", x"10", x"32", x"7F", x"7E", x"3C", x"38", x"3E", x"34", x"1E", x"1E", x"34", x"2C", x"08", x"00", x"3E", x"34", x"1E", x"1E", x"04", x"40", x"40", x"0C", x"0C", x"1E", x"1C", x"0C", x"00", x"81", x"C3", x"42", x"0C", x"1E", x"10", x"32", x"7F", x"7E", x"3C", x"3C", x"3C", x"3C", x"1C", x"18", x"08", x"08", x"10", x"00", x"3C", x"3C", x"1C", x"08", x"10", x"10", x"20", x"10", x"0C", x"1E", x"1C", x"0C", x"00", x"C1", x"61", x"32", x"0C", x"1E", x"10", x"32", x"7F", x"3E", x"1E", x"0C", x"3C", x"3C", x"36", x"66", x"66", x"46", x"02", x"00", x"3C", x"3C", x"36", x"66", x"24", x"80", x"84", x"03", x"00", x"0C", x"1E", x"04", x"00", x"00", x"19", x"0E", x"00", x"0C", x"1E", x"38", x"3C", x"7C", x"60", x"70", 
															x"38", x"38", x"1C", x"3C", x"7C", x"58", x"08", x"00", x"38", x"38", x"1C", x"3C", x"1C", x"80", x"50", x"0C", x"1C", x"1E", x"1F", x"3B", x"33", x"63", x"42", x"00", x"1C", x"1E", x"1F", x"3B", x"12", x"00", x"80", x"63", x"01", x"03", x"1D", x"3D", x"00", x"80", x"C0", x"40", x"00", x"00", x"1C", x"3A", x"7F", x"7E", x"3C", x"3C", x"01", x"03", x"1D", x"3D", x"00", x"80", x"80", x"00", x"00", x"00", x"1C", x"3A", x"7F", x"7E", x"3C", x"3C", x"01", x"03", x"19", x"3D", x"00", x"80", x"C0", x"40", x"00", x"00", x"18", x"3E", x"7F", x"7E", x"3C", x"3C", x"01", x"03", x"19", x"3D", x"00", x"80", x"80", x"00", x"00", x"00", x"18", x"3E", x"7F", x"7E", x"3C", x"3C", x"01", x"1B", x"3D", x"39", x"19", x"00", x"80", x"60", x"00", x"18", x"3C", x"20", x"66", x"FE", x"7C", x"1C", x"01", x"1B", x"3D", x"39", x"19", x"00", x"80", x"80", x"00", x"18", x"3C", x"20", x"66", x"FE", x"7C", x"7C", 
															x"01", x"1B", x"3D", x"3D", x"19", x"00", x"80", x"60", x"00", x"18", x"3C", x"24", x"66", x"FE", x"7C", x"1C", x"01", x"1B", x"3D", x"3D", x"19", x"00", x"80", x"80", x"00", x"18", x"3C", x"24", x"66", x"FE", x"7C", x"7C", x"00", x"00", x"00", x"18", x"3C", x"00", x"80", x"C2", x"00", x"00", x"00", x"18", x"3C", x"7E", x"7F", x"3C", x"00", x"00", x"18", x"3C", x"3C", x"18", x"81", x"63", x"00", x"00", x"18", x"3C", x"66", x"E7", x"7E", x"1C", x"18", x"3C", x"1C", x"18", x"00", x"81", x"81", x"C3", x"18", x"3C", x"04", x"66", x"FF", x"3C", x"3C", x"3C", x"00", x"18", x"3C", x"00", x"00", x"00", x"C1", x"03", x"00", x"18", x"3C", x"7C", x"FE", x"FF", x"3C", x"3C", x"F8", x"F8", x"6C", x"3C", x"6C", x"46", x"40", x"00", x"F8", x"F8", x"6C", x"3C", x"00", x"80", x"83", x"40", x"F8", x"D8", x"7C", x"3E", x"36", x"62", x"00", x"00", x"F8", x"D8", x"7C", x"3E", x"00", x"00", x"C3", x"00", 
															x"00", x"00", x"00", x"18", x"3C", x"00", x"C3", x"42", x"00", x"00", x"00", x"18", x"3C", x"7E", x"3C", x"3C", x"7C", x"EC", x"C6", x"46", x"02", x"00", x"00", x"00", x"7C", x"EC", x"06", x"04", x"C1", x"02", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"99", x"81", x"42", x"00", x"00", x"18", x"3C", x"66", x"66", x"7E", x"3C", x"3C", x"6E", x"C6", x"66", x"24", x"00", x"00", x"00", x"3C", x"6E", x"C6", x"0E", x"08", x"64", x"00", x"00", x"00", x"0C", x"1E", x"1C", x"0C", x"80", x"C1", x"63", x"00", x"0C", x"1E", x"30", x"72", x"7F", x"3E", x"1C", x"3C", x"36", x"1B", x"1B", x"36", x"20", x"00", x"00", x"3C", x"36", x"1B", x"1B", x"00", x"44", x"22", x"00", x"00", x"00", x"18", x"3C", x"00", x"20", x"61", x"C0", x"00", x"00", x"18", x"3C", x"3E", x"1F", x"1E", x"1E", x"1E", x"36", x"6C", x"66", x"22", x"00", x"00", x"00", x"1E", x"36", x"6C", x"00", x"11", x"66", x"00", x"00", 
															x"00", x"00", x"30", x"78", x"38", x"00", x"90", x"F0", x"00", x"00", x"30", x"78", x"18", x"3C", x"2E", x"0E", x"1E", x"36", x"6C", x"6C", x"36", x"12", x"00", x"00", x"1E", x"36", x"6C", x"6C", x"00", x"01", x"36", x"00", x"00", x"00", x"00", x"18", x"3C", x"00", x"01", x"81", x"00", x"00", x"00", x"18", x"3C", x"7E", x"FE", x"7C", x"F8", x"6C", x"6C", x"64", x"40", x"00", x"00", x"00", x"F8", x"6C", x"6C", x"20", x"86", x"80", x"00", x"00", x"00", x"00", x"60", x"F0", x"60", x"00", x"90", x"70", x"00", x"00", x"60", x"F0", x"38", x"7C", x"6E", x"0E", x"3E", x"7E", x"6C", x"26", x"00", x"00", x"00", x"00", x"3E", x"7E", x"0C", x"01", x"61", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"00", x"01", x"41", x"C0", x"00", x"00", x"18", x"3C", x"3E", x"7E", x"3E", x"3E", x"7C", x"F8", x"6E", x"0C", x"00", x"00", x"00", x"00", x"7C", x"FA", x"09", x"E9", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"18", x"3C", x"3C", x"98", x"81", x"C1", x"00", x"00", x"18", x"3C", x"66", x"67", x"3C", x"3C", x"3C", x"6C", x"6C", x"24", x"00", x"00", x"00", x"00", x"3C", x"6C", x"0C", x"02", x"62", x"00", x"00", x"00", x"00", x"18", x"3C", x"1C", x"18", x"00", x"62", x"CE", x"00", x"18", x"3C", x"04", x"26", x"3F", x"1D", x"10", x"3E", x"6C", x"36", x"10", x"00", x"00", x"00", x"00", x"3E", x"6C", x"21", x"09", x"30", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"0C", x"7E", x"FF", x"FF", x"00", x"00", x"00", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"7E", x"FF", x"FF", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"81", x"C3", x"66", x"18", x"3C", x"24", x"66", x"FF", x"7E", x"3C", x"18", 
															x"3E", x"36", x"36", x"63", x"63", x"63", x"22", x"00", x"3E", x"36", x"36", x"63", x"22", x"00", x"00", x"63", x"0C", x"1E", x"1C", x"00", x"01", x"0B", x"0E", x"00", x"0C", x"1E", x"18", x"3C", x"7C", x"74", x"70", x"3C", x"0C", x"1E", x"1C", x"00", x"00", x"01", x"2C", x"38", x"0C", x"1E", x"18", x"3C", x"7E", x"7E", x"52", x"04", x"0C", x"1E", x"1C", x"00", x"01", x"83", x"C0", x"60", x"0C", x"1E", x"18", x"3C", x"7C", x"7C", x"3C", x"1C", x"3C", x"3E", x"1F", x"3B", x"32", x"62", x"40", x"00", x"3C", x"3E", x"1F", x"3A", x"30", x"04", x"83", x"60", x"3C", x"38", x"1C", x"3C", x"3C", x"2C", x"24", x"00", x"3C", x"38", x"1C", x"1C", x"08", x"40", x"40", x"26", x"3C", x"3C", x"1E", x"36", x"76", x"02", x"02", x"00", x"3C", x"3C", x"1E", x"36", x"94", x"80", x"00", x"03", x"06", x"1B", x"FD", x"BD", x"81", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"7E", x"FF", x"7E", x"3C", 
															x"66", x"DB", x"BD", x"BD", x"18", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"FF", x"FF", x"7E", x"3C", x"3C", x"3E", x"36", x"36", x"34", x"24", x"00", x"00", x"3C", x"3E", x"36", x"36", x"58", x"48", x"48", x"00", x"3E", x"77", x"63", x"63", x"63", x"22", x"00", x"00", x"3E", x"77", x"63", x"00", x"00", x"00", x"63", x"00", x"00", x"00", x"18", x"3C", x"00", x"81", x"C3", x"00", x"00", x"00", x"18", x"3C", x"7E", x"7E", x"3C", x"3C", x"7C", x"6C", x"36", x"36", x"32", x"20", x"00", x"00", x"7C", x"6C", x"36", x"34", x"04", x"44", x"30", x"00", x"00", x"00", x"18", x"3C", x"00", x"81", x"81", x"C3", x"00", x"00", x"18", x"3C", x"7E", x"7E", x"34", x"3C", x"3C", x"7E", x"76", x"32", x"30", x"20", x"20", x"00", x"3C", x"7E", x"75", x"31", x"00", x"00", x"00", x"30", x"3C", x"7E", x"E7", x"C3", x"C3", x"42", x"00", x"00", x"FF", x"FF", x"E7", x"C3", x"00", x"00", x"C3", x"00", 
															x"3C", x"76", x"66", x"63", x"07", x"06", x"04", x"00", x"3C", x"76", x"66", x"A3", x"43", x"40", x"00", x"06", x"00", x"18", x"3C", x"3C", x"18", x"81", x"87", x"CC", x"00", x"18", x"3C", x"66", x"E7", x"7E", x"78", x"30", x"5C", x"5E", x"16", x"06", x"06", x"04", x"04", x"00", x"7C", x"7E", x"36", x"06", x"04", x"00", x"00", x"06", x"C6", x"B2", x"FA", x"BA", x"32", x"00", x"00", x"00", x"00", x"30", x"78", x"18", x"CC", x"7E", x"7C", x"3C", x"3C", x"7C", x"68", x"78", x"3C", x"16", x"02", x"00", x"3C", x"7C", x"68", x"18", x"00", x"00", x"31", x"06", x"18", x"3C", x"1C", x"18", x"40", x"40", x"2C", x"18", x"18", x"3C", x"0C", x"24", x"3E", x"3E", x"12", x"06", x"1E", x"1E", x"34", x"34", x"1A", x"0E", x"00", x"00", x"1E", x"1E", x"34", x"34", x"00", x"01", x"05", x"04", x"00", x"18", x"3C", x"1C", x"18", x"00", x"40", x"38", x"00", x"18", x"3C", x"0C", x"04", x"3E", x"3E", x"06", 
															x"0E", x"1E", x"3C", x"2C", x"36", x"12", x"12", x"00", x"0E", x"1E", x"3C", x"2C", x"00", x"00", x"01", x"36", x"43", x"99", x"BD", x"9D", x"18", x"00", x"00", x"00", x"00", x"18", x"3C", x"04", x"E7", x"7E", x"3C", x"3C", x"3C", x"3C", x"6C", x"78", x"5C", x"6C", x"24", x"00", x"3C", x"3C", x"6C", x"78", x"18", x"00", x"02", x"64", x"00", x"00", x"00", x"00", x"66", x"66", x"76", x"7E", x"00", x"00", x"00", x"66", x"00", x"24", x"76", x"7E", x"3E", x"7E", x"EC", x"D8", x"4C", x"64", x"20", x"00", x"3E", x"7E", x"EC", x"D8", x"00", x"02", x"12", x"24", x"00", x"00", x"18", x"3C", x"3C", x"18", x"82", x"F6", x"00", x"00", x"18", x"3C", x"66", x"E7", x"7D", x"08", x"7E", x"E7", x"C3", x"C3", x"42", x"00", x"00", x"00", x"7E", x"E7", x"C3", x"00", x"00", x"C3", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"7E", x"FF", x"FF", 
															x"3C", x"7E", x"E7", x"C3", x"C3", x"42", x"00", x"00", x"FF", x"7F", x"E7", x"F3", x"00", x"00", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"78", x"78", x"00", x"00", x"00", x"00", x"00", x"30", x"7E", x"CF", x"FF", x"BF", x"0E", x"00", x"00", x"81", x"81", x"3C", x"18", x"7C", x"FC", x"FE", x"FF", x"7E", x"7E", x"00", x"3E", x"7E", x"E7", x"C3", x"43", x"02", x"00", x"00", x"3E", x"7E", x"E7", x"03", x"00", x"C0", x"03", x"00", x"0C", x"1E", x"5E", x"4C", x"60", x"01", x"01", x"00", x"0C", x"1E", x"1E", x"0C", x"1F", x"3E", x"1E", x"1E", x"1C", x"18", x"30", x"30", x"10", x"10", x"00", x"00", x"1C", x"18", x"30", x"00", x"60", x"00", x"30", x"00", x"40", x"4C", x"7E", x"3E", x"0C", x"00", x"01", x"06", x"00", x"0C", x"1E", x"1E", x"3E", x"1F", x"1E", x"18", x"1E", x"34", x"6C", x"66", x"62", x"20", x"00", x"00", x"1E", x"34", x"6C", x"00", x"00", x"06", x"60", x"00", 
															x"98", x"BC", x"F8", x"40", x"00", x"00", x"03", x"00", x"18", x"3C", x"30", x"38", x"3C", x"7C", x"7C", x"3C", x"00", x"18", x"3C", x"39", x"03", x"0E", x"80", x"00", x"00", x"18", x"3C", x"30", x"78", x"F0", x"78", x"78", x"3C", x"7E", x"E7", x"C3", x"C3", x"42", x"00", x"00", x"FF", x"7E", x"E7", x"E7", x"00", x"00", x"C3", x"00", x"00", x"00", x"00", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"7E", x"FF", x"FF", x"3C", x"7E", x"E7", x"C3", x"C3", x"42", x"00", x"00", x"FF", x"7E", x"E7", x"E7", x"24", x"00", x"C3", x"00", x"18", x"3C", x"BD", x"99", x"81", x"C3", x"00", x"00", x"7E", x"FF", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"18", x"4C", x"66", x"3C", x"18", x"00", x"30", x"00", x"C0", x"0C", x"06", x"3C", x"18", x"00", x"00", x"00", x"0C", x"1E", x"1C", x"0C", x"21", x"3B", x"00", x"30", x"7C", x"FE", x"73", x"33", x"00", x"00", 
															x"00", x"00", x"07", x"7F", x"37", x"1C", x"30", x"00", x"00", x"00", x"07", x"9F", x"97", x"0C", x"40", x"40", x"18", x"3E", x"18", x"01", x"07", x"00", x"00", x"00", x"18", x"3C", x"F0", x"F8", x"F8", x"18", x"00", x"00", x"04", x"0E", x"1B", x"37", x"6E", x"1C", x"10", x"00", x"04", x"0E", x"1B", x"17", x"8E", x"84", x"20", x"20", x"0C", x"1D", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"2C", x"3E", x"7C", x"FC", x"F0", x"60", x"00", x"00", x"00", x"66", x"DB", x"BD", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"FF", x"7E", x"7E", x"3E", x"7E", x"E7", x"C3", x"66", x"24", x"00", x"00", x"3E", x"7E", x"E7", x"C3", x"00", x"08", x"66", x"00", x"18", x"38", x"18", x"38", x"2A", x"AA", x"AB", x"AE", x"18", x"38", x"00", x"24", x"7E", x"FF", x"3C", x"38", x"3C", x"7C", x"EC", x"CC", x"C6", x"63", x"21", x"60", x"3C", x"7C", x"EC", x"CC", x"02", x"62", x"20", x"00", 
															x"18", x"38", x"18", x"38", x"2A", x"AA", x"E9", x"6B", x"18", x"38", x"00", x"24", x"7E", x"7F", x"3C", x"3C", x"1C", x"1C", x"3C", x"38", x"18", x"18", x"0C", x"18", x"1C", x"1C", x"3C", x"38", x"00", x"18", x"08", x"00", x"18", x"38", x"18", x"38", x"AA", x"AA", x"A9", x"EB", x"18", x"38", x"00", x"24", x"FE", x"FF", x"7C", x"1C", x"3C", x"3C", x"18", x"38", x"3C", x"36", x"24", x"60", x"3C", x"3C", x"18", x"38", x"0C", x"34", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"98", x"B8", x"98", x"38", x"2A", x"2B", x"29", x"2B", x"18", x"38", x"40", x"64", x"3F", x"3E", x"3C", x"3C", x"1C", x"1C", x"14", x"14", x"14", x"14", x"36", x"00", x"1C", x"1C", x"14", x"00", x"14", x"14", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"81", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"99", x"B9", x"9B", x"3A", x"28", x"28", x"28", x"28", x"18", x"38", x"42", x"66", x"3C", x"3C", x"3C", x"3C", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"B8", x"2A", x"2A", x"2A", x"2E", x"18", x"38", x"00", x"64", x"7E", x"3E", x"3C", x"30", x"3C", x"38", x"38", x"38", x"28", x"28", x"78", x"00", x"3C", x"38", x"38", x"00", x"28", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"00", x"00", x"38", x"10", x"38", x"7C", x"FE", x"FE", x"38", x"38", x"38", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"08", x"00", x"00", x"00", x"08", x"1C", x"1C", x"1C", x"1C", x"08", x"00", x"00", x"00", x"1C", x"00", x"00", x"1C", x"00", x"00", x"08", x"1C", x"3E", x"3E", x"3E", x"3E", x"1C", x"08", 
															x"00", x"00", x"00", x"00", x"00", x"1C", x"00", x"00", x"00", x"00", x"00", x"08", x"1C", x"3E", x"3E", x"3E", x"00", x"00", x"00", x"22", x"36", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"00", x"00", x"00", x"00", x"00", x"3E", x"3E", x"3E", x"1C", x"08", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"81", x"E1", x"32", x"18", x"3C", x"24", x"66", x"FF", x"7E", x"1E", x"0C", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"7E", x"3C", x"00", x"00", x"30", x"78", x"00", x"00", x"01", x"01", x"C0", x"00", x"30", x"78", x"7C", x"FE", x"7E", x"7E", x"3E", x"00", x"30", x"78", x"00", x"00", x"00", x"01", x"60", x"00", x"30", x"78", x"7C", x"FE", x"FF", x"7E", x"1E", 
															x"00", x"30", x"78", x"00", x"00", x"00", x"32", x"60", x"00", x"30", x"78", x"7C", x"FE", x"7E", x"0C", x"1C", x"0F", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"F0", x"F8", x"FC", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0E", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"80", x"00", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"F0", x"70", x"30", x"10", x"FF", x"7F", x"3F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"08", x"0C", x"0E", x"0F", x"0F", x"0F", x"0F", 
															x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0E", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"07", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0F", x"F8", x"FC", x"FE", x"FF", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"FF", x"F7", x"F3", x"F1", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0E", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"1F", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"00", x"80", x"C0", x"E0", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F8", x"FC", x"FE", x"0F", x"0F", x"0F", x"0F", x"0F", x"07", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"1F", x"F8", x"70", x"38", x"1C", x"1C", x"0E", x"07", x"07", x"F8", x"70", x"38", x"1C", x"1C", x"0E", x"07", x"07", x"0F", x"07", x"0E", x"1C", x"1C", x"38", x"70", x"70", x"0F", x"07", x"0E", x"1C", x"1C", x"38", x"70", x"70", x"9C", x"1C", x"3E", x"36", x"77", x"77", x"E3", x"E3", x"9C", x"1C", x"3E", x"36", x"77", x"77", x"E3", x"E3", x"07", x"03", x"03", x"03", x"03", x"03", x"83", x"83", x"07", x"03", x"03", x"03", x"03", x"03", x"83", x"83", x"FE", x"FF", x"83", x"81", x"81", x"81", x"83", x"FF", x"FE", x"FF", x"83", x"81", x"81", x"81", x"83", x"FF", 
															x"1F", x"0F", x"8E", x"CE", x"CE", x"CE", x"8E", x"0E", x"1F", x"0F", x"8E", x"CE", x"CE", x"CE", x"8E", x"0E", x"F0", x"F8", x"1C", x"0C", x"0E", x"0E", x"0E", x"0E", x"F0", x"F8", x"1C", x"0C", x"0E", x"0E", x"0E", x"0E", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"E0", x"C1", x"C1", x"C1", x"C3", x"C3", x"C3", x"E7", x"E0", x"C1", x"C1", x"C1", x"C3", x"C3", x"C3", x"E7", x"E3", x"C1", x"FF", x"FF", x"80", x"80", x"80", x"C1", x"E3", x"C1", x"FF", x"FF", x"80", x"80", x"80", x"C1", x"83", x"C3", x"C3", x"C3", x"E3", x"E3", x"E3", x"F7", x"83", x"C3", x"C3", x"C3", x"E3", x"E3", x"E3", x"F7", x"FE", x"87", x"83", x"83", x"83", x"83", x"83", x"C3", x"FE", x"87", x"83", x"83", x"83", x"83", x"83", x"C3", x"0E", x"0E", x"8E", x"8E", x"8E", x"8E", x"8F", x"DF", x"0E", x"0E", x"8E", x"8E", x"8E", x"8E", x"8F", x"DF", 
															x"00", x"0E", x"08", x"08", x"0E", x"02", x"02", x"0E", x"00", x"0E", x"08", x"08", x"0E", x"02", x"02", x"0E", x"00", x"EE", x"AA", x"AA", x"AA", x"AA", x"AA", x"EE", x"00", x"EE", x"AA", x"AA", x"AA", x"AA", x"AA", x"EE", x"00", x"EE", x"8A", x"8A", x"EA", x"2A", x"2A", x"EE", x"00", x"EE", x"8A", x"8A", x"EA", x"2A", x"2A", x"EE", x"00", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"00", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"00", x"0C", x"12", x"02", x"02", x"04", x"08", x"1E", x"00", x"0C", x"12", x"02", x"02", x"04", x"08", x"1E", x"00", x"4E", x"48", x"48", x"4E", x"42", x"42", x"4E", x"00", x"4E", x"48", x"48", x"4E", x"42", x"42", x"4E", x"0E", x"0E", x"0E", x"0E", x"0C", x"1C", x"F8", x"F0", x"0E", x"0E", x"0E", x"0E", x"0C", x"1C", x"F8", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00", x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00", x"0C", x"1C", x"0C", x"0C", x"0C", x"0C", x"3F", x"00", x"0C", x"1C", x"0C", x"0C", x"0C", x"0C", x"3F", x"00", x"3E", x"63", x"07", x"1E", x"3C", x"70", x"7F", x"00", x"3E", x"63", x"07", x"1E", x"3C", x"70", x"7F", x"00", x"3F", x"06", x"0C", x"1E", x"03", x"63", x"3E", x"00", x"3F", x"06", x"0C", x"1E", x"03", x"63", x"3E", x"00", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"7E", x"60", x"7E", x"03", x"03", x"63", x"3E", x"00", x"7E", x"60", x"7E", x"03", x"03", x"63", x"3E", x"00", x"1E", x"30", x"60", x"7E", x"63", x"63", x"3E", x"00", x"1E", x"30", x"60", x"7E", x"63", x"63", x"3E", x"00", x"7F", x"63", x"06", x"0C", x"18", x"18", x"18", x"00", x"7F", x"63", x"06", x"0C", x"18", x"18", x"18", x"00", 
															x"3C", x"62", x"72", x"3C", x"4F", x"43", x"3E", x"00", x"3C", x"62", x"72", x"3C", x"4F", x"43", x"3E", x"00", x"3E", x"63", x"63", x"3F", x"03", x"06", x"3C", x"00", x"3E", x"63", x"63", x"3F", x"03", x"06", x"3C", x"00", x"1C", x"36", x"63", x"63", x"7F", x"63", x"63", x"00", x"1C", x"36", x"63", x"63", x"7F", x"63", x"63", x"00", x"7E", x"63", x"63", x"7E", x"63", x"63", x"7E", x"00", x"7E", x"63", x"63", x"7E", x"63", x"63", x"7E", x"00", x"1E", x"33", x"60", x"60", x"60", x"33", x"1E", x"00", x"1E", x"33", x"60", x"60", x"60", x"33", x"1E", x"00", x"7C", x"66", x"63", x"63", x"63", x"66", x"7C", x"00", x"7C", x"66", x"63", x"63", x"63", x"66", x"7C", x"00", x"3F", x"30", x"30", x"3E", x"30", x"30", x"3F", x"00", x"3F", x"30", x"30", x"3E", x"30", x"30", x"3F", x"00", x"7F", x"60", x"60", x"7E", x"60", x"60", x"60", x"00", x"7F", x"60", x"60", x"7E", x"60", x"60", x"60", x"00", 
															x"1F", x"30", x"60", x"67", x"63", x"33", x"1F", x"00", x"1F", x"30", x"60", x"67", x"63", x"33", x"1F", x"00", x"63", x"63", x"63", x"7F", x"63", x"63", x"63", x"00", x"63", x"63", x"63", x"7F", x"63", x"63", x"63", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"0C", x"1E", x"00", x"03", x"03", x"03", x"03", x"03", x"63", x"3E", x"00", x"03", x"03", x"03", x"03", x"03", x"63", x"3E", x"00", x"63", x"66", x"6C", x"78", x"7C", x"6E", x"67", x"00", x"63", x"66", x"6C", x"78", x"7C", x"6E", x"67", x"00", x"30", x"30", x"30", x"30", x"30", x"30", x"3F", x"00", x"30", x"30", x"30", x"30", x"30", x"30", x"3F", x"00", x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00", x"63", x"77", x"7F", x"7F", x"6B", x"63", x"63", x"00", x"63", x"73", x"7B", x"7F", x"6F", x"67", x"63", x"00", x"63", x"73", x"7B", x"7F", x"6F", x"67", x"63", x"00", 
															x"3E", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"3E", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"7E", x"63", x"63", x"63", x"7E", x"60", x"60", x"00", x"7E", x"63", x"63", x"63", x"7E", x"60", x"60", x"00", x"3E", x"63", x"63", x"63", x"6F", x"66", x"3D", x"00", x"3E", x"63", x"63", x"63", x"6F", x"66", x"3D", x"00", x"7E", x"63", x"63", x"67", x"7C", x"6E", x"67", x"00", x"7E", x"63", x"63", x"67", x"7C", x"6E", x"67", x"00", x"3C", x"66", x"60", x"3E", x"03", x"63", x"3E", x"00", x"3C", x"66", x"60", x"3E", x"03", x"63", x"3E", x"00", x"3F", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"3F", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"63", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"63", x"63", x"63", x"63", x"63", x"63", x"3E", x"00", x"63", x"63", x"63", x"77", x"3E", x"1C", x"08", x"00", x"63", x"63", x"63", x"77", x"3E", x"1C", x"08", x"00", 
															x"63", x"63", x"6B", x"7F", x"7F", x"36", x"22", x"00", x"63", x"63", x"6B", x"7F", x"7F", x"36", x"22", x"00", x"63", x"77", x"3E", x"1C", x"3E", x"77", x"63", x"00", x"63", x"77", x"3E", x"1C", x"3E", x"77", x"63", x"00", x"33", x"33", x"12", x"1E", x"0C", x"0C", x"0C", x"00", x"33", x"33", x"12", x"1E", x"0C", x"0C", x"0C", x"00", x"7F", x"07", x"0E", x"1C", x"38", x"70", x"7F", x"00", x"7F", x"07", x"0E", x"1C", x"38", x"70", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"7E", x"00", x"00", x"7E", x"00", x"00", x"00", x"00", x"7E", x"00", x"00", x"7E", x"00", x"00", x"6C", x"6C", x"6C", x"6C", x"00", x"6C", x"6C", x"00", x"6C", x"6C", x"6C", x"6C", x"00", x"6C", x"6C", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"08", x"18", x"5A", x"3C", x"18", x"3C", x"5A", x"18", x"00", x"18", x"5A", x"3C", x"18", x"3C", x"5A", x"18", x"00", x"0C", x"18", x"30", x"60", x"30", x"18", x"0C", x"00", x"0C", x"18", x"30", x"60", x"30", x"18", x"0C", x"00", x"30", x"18", x"0C", x"06", x"0C", x"18", x"30", x"00", x"30", x"18", x"0C", x"06", x"0C", x"18", x"30", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"67", x"6C", x"2C", x"47", x"00", x"08", x"07", x"00", x"67", x"6C", x"2C", x"47", x"00", x"08", x"07", x"00", x"80", x"C0", x"00", x"80", x"C0", x"C0", x"80", x"00", x"80", x"C0", x"00", x"80", x"C0", x"C0", x"80", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"7E", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", x"81", x"81", x"81", x"81", x"FF", x"81", x"81", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"81", x"81", x"81", x"81", x"81", x"81", x"81", 
															x"00", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"7E", x"7E", x"7E", x"00", x"7E", x"7E", x"7E", x"81", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"7E", x"7E", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"81", x"81", x"81", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"81", x"81", x"81", x"81", x"FF", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1C", x"30", x"60", x"C1", x"83", x"07", x"00", x"00", x"03", x"0F", x"1F", x"3E", x"7C", x"F8", x"FF", x"80", x"00", x"00", x"7F", x"FF", x"FF", x"80", x"00", x"7F", x"FF", x"FF", x"80", x"00", x"00", x"00", x"80", x"F0", x"1C", x"06", x"03", x"C1", x"E0", x"F0", x"00", x"00", x"E0", x"F8", x"FC", x"3E", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"02", x"06", x"04", x"04", x"0C", x"08", x"08", x"18", x"01", x"01", x"03", x"03", x"03", x"07", x"07", x"07", x"0F", x"1C", x"38", x"38", x"70", x"70", x"E0", x"E0", x"F0", x"E0", x"C0", x"C0", x"80", x"80", x"00", x"00", x"78", x"1C", x"0E", x"0E", x"07", x"07", x"03", x"03", x"07", x"03", x"01", x"01", x"00", x"00", x"00", x"00", 
															x"20", x"30", x"10", x"10", x"18", x"08", x"88", x"88", x"C0", x"C0", x"E0", x"E0", x"E0", x"F0", x"70", x"70", x"11", x"11", x"1F", x"00", x"00", x"00", x"00", x"00", x"0E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"E0", x"38", x"0C", x"04", x"06", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"03", x"03", x"03", x"03", x"83", x"43", x"43", x"83", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"8C", x"84", x"84", x"84", x"84", x"8C", x"88", x"88", x"70", x"78", x"78", x"78", x"78", x"70", x"70", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"02", x"02", x"02", x"00", x"00", x"03", x"1D", x"E0", x"00", x"00", x"00", x"03", x"1F", x"FC", x"E0", x"01", 
															x"00", x"00", x"00", x"10", x"28", x"14", x"08", x"30", x"00", x"00", x"70", x"E8", x"D4", x"68", x"F0", x"C0", x"03", x"03", x"03", x"03", x"03", x"07", x"0C", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"88", x"88", x"B8", x"E0", x"80", x"00", x"00", x"00", x"70", x"70", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"01", x"00", x"00", x"00", x"00", x"01", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"07", x"38", x"C4", x"02", x"01", x"00", x"00", x"00", x"F8", x"C7", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"04", x"88", x"10", x"60", x"03", x"07", x"8E", x"DC", x"F8", x"70", x"E0", x"00", x"40", x"E0", x"31", x"1F", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"8C", x"07", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"06", x"08", x"11", x"20", x"40", x"80", x"00", x"00", x"00", x"07", x"0E", x"1F", x"3B", x"71", x"E0", x"C0", x"00", x"00", x"00", x"80", x"40", x"23", x"1C", x"E0", x"00", x"00", x"00", x"00", x"80", x"C0", x"E3", x"1F", x"00", x"00", x"00", x"00", x"80", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"80", x"00", x"00", x"00", x"01", x"07", x"1D", x"11", x"11", x"00", x"00", x"00", x"00", x"00", x"02", x"0E", x"0E", x"18", x"30", x"60", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"10", x"28", x"14", x"08", x"00", x"00", x"00", x"03", x"0F", x"16", x"2B", x"17", x"0E", x"00", x"00", 
															x"07", x"B8", x"C0", x"00", x"00", x"40", x"40", x"40", x"80", x"07", x"3F", x"F8", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"11", x"11", x"31", x"21", x"21", x"21", x"21", x"31", x"0E", x"0E", x"0E", x"1E", x"1E", x"1E", x"1E", x"0E", x"C1", x"C2", x"C2", x"C1", x"C0", x"C0", x"C0", x"C0", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"80", x"40", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"40", x"60", x"20", x"30", x"1C", x"07", x"07", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"88", x"88", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"70", x"10", x"10", x"10", x"18", x"08", x"08", x"0C", x"04", x"0F", x"0F", x"0F", x"07", x"07", x"07", x"03", x"03", 
															x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"01", x"08", x"08", x"1C", x"1C", x"3E", x"FF", x"FF", x"FF", x"08", x"08", x"1C", x"1C", x"3E", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"02", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"02", x"FF", x"FF", x"FF", x"F7", x"E3", x"80", x"00", x"00", x"FF", x"FF", x"FF", x"F7", x"E3", x"80", x"00", x"00", x"80", x"80", x"80", x"C0", x"C0", x"E0", x"60", x"20", x"80", x"80", x"80", x"C0", x"C0", x"E0", x"60", x"20", x"00", x"00", x"00", x"00", x"08", x"08", x"1C", x"1C", x"08", x"08", x"08", x"1C", x"1C", x"3E", x"3E", x"7F", x"00", x"0F", x"07", x"01", x"00", x"00", x"00", x"01", x"7F", x"3F", x"1F", x"0F", x"03", x"01", x"03", x"03", 
															x"3E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"02", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07", x"0F", x"0C", x"18", x"10", x"00", x"F8", x"F0", x"C0", x"80", x"80", x"80", x"C0", x"FF", x"FE", x"FC", x"F8", x"E0", x"C0", x"E0", x"E0", x"E3", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"F7", x"E3", x"80", x"00", x"00", x"00", x"00", x"C0", x"E0", x"60", x"20", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"78", x"18", x"0C", x"04", x"04", x"04", x"06", x"07", x"0F", x"1F", x"3F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"F8", x"FE", x"FF", x"00", x"10", x"28", x"1A", x"0D", x"06", x"01", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1C", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"3F", x"7F", x"3F", x"3E", x"18", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"80", x"80", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"0C", x"07", x"07", x"07", x"1C", x"38", x"80", x"C6", x"F3", x"00", x"00", x"00", x"00", x"00", 
															x"78", x"70", x"E0", x"E0", x"80", x"F8", x"F8", x"18", x"03", x"03", x"06", x"0C", x"18", x"00", x"00", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0D", x"07", x"07", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"F8", x"02", x"06", x"0E", x"1C", x"38", x"74", x"FC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"7C", x"FF", x"9F", x"37", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"0F", x"0F", x"1F", x"3F", x"FF", x"FF", x"F8", x"F8", x"F0", x"F0", x"60", x"00", x"00", x"00", x"F4", x"F8", x"F0", x"F0", x"E0", x"C0", x"86", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"07", x"05", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"0D", x"01", x"02", x"FF", x"FF", x"FF", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"88", x"3C", x"64", x"FE", x"F8", x"F4", x"F8", x"D0", x"60", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"18", x"3F", x"3F", x"3F", x"17", x"38", x"7C", x"FE", x"FC", x"E0", x"00", x"00", x"03", x"00", x"00", x"00", x"03", x"1F", x"FF", x"FF", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FE", x"7E", x"03", x"01", x"00", x"00", x"07", x"07", x"0F", x"0C", x"0C", x"0E", x"07", x"07", x"00", x"00", x"00", x"03", x"F8", x"E1", x"03", x"87", x"8F", x"DF", x"FF", x"3F", x"07", x"1E", x"FC", x"78", x"70", x"20", x"00", x"C0", 
															x"00", x"60", x"F0", x"F0", x"E0", x"C0", x"80", x"00", x"FC", x"98", x"00", x"00", x"00", x"04", x"0C", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"00", x"00", x"01", x"03", x"1F", x"07", x"9E", x"FC", x"EC", x"0C", x"1C", x"00", x"00", x"00", x"60", x"00", x"13", x"F3", x"E3", x"FE", x"FC", x"F0", x"00", x"00", x"40", x"40", x"00", x"00", x"00", x"00", x"18", x"30", x"B0", x"9C", x"0E", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BB", x"BB", x"BB", x"1B", x"B9", x"BA", x"BA", x"CA", x"44", x"44", x"44", x"E4", x"46", x"45", x"45", x"35", 
															x"FF", x"FF", x"FF", x"FF", x"BB", x"BB", x"BB", x"1B", x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"E4", x"B9", x"BA", x"BA", x"CA", x"FF", x"FF", x"FF", x"FF", x"46", x"45", x"45", x"35", x"00", x"00", x"00", x"00", x"FB", x"FB", x"FB", x"90", x"7B", x"9B", x"EB", x"1C", x"04", x"04", x"04", x"6F", x"84", x"64", x"14", x"E3", x"FE", x"FE", x"FE", x"B8", x"56", x"56", x"56", x"58", x"01", x"01", x"01", x"47", x"A9", x"A9", x"A9", x"A7", x"FE", x"FE", x"FE", x"58", x"36", x"76", x"76", x"78", x"01", x"01", x"01", x"A7", x"C9", x"89", x"89", x"87", x"CF", x"B7", x"B6", x"CD", x"B3", x"7B", x"75", x"8E", x"30", x"48", x"49", x"32", x"4C", x"84", x"8A", x"71", x"FF", x"E7", x"E7", x"FF", x"E7", x"E7", x"FF", x"FF", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"90", x"00", x"00", x"00", x"00", x"04", x"04", x"04", x"6F", 
															x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"B8", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"47", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"58", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"A7", x"FF", x"FF", x"FF", x"FF", x"CF", x"B7", x"B6", x"CD", x"00", x"00", x"00", x"00", x"30", x"48", x"49", x"32", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"FF", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"7B", x"9B", x"EB", x"1C", x"FF", x"FF", x"FF", x"FF", x"84", x"64", x"14", x"E3", x"00", x"00", x"00", x"00", x"56", x"56", x"56", x"58", x"FF", x"FF", x"FF", x"FF", x"A9", x"A9", x"A9", x"A7", x"00", x"00", x"00", x"00", x"36", x"76", x"76", x"78", x"FF", x"FF", x"FF", x"FF", x"C9", x"89", x"89", x"87", x"00", x"00", x"00", x"00", x"B3", x"7B", x"75", x"8E", x"FF", x"FF", x"FF", x"FF", x"4C", x"84", x"8A", x"71", x"00", x"00", x"00", x"00", 
															x"E7", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"E3", x"C9", x"9C", x"9C", x"9C", x"C9", x"E3", x"FF", x"1C", x"36", x"63", x"63", x"63", x"36", x"1C", x"00", x"F3", x"E3", x"F3", x"F3", x"F3", x"F3", x"C0", x"FF", x"0C", x"1C", x"0C", x"0C", x"0C", x"0C", x"3F", x"00", x"C1", x"9C", x"F8", x"E1", x"C3", x"8F", x"80", x"FF", x"3E", x"63", x"07", x"1E", x"3C", x"70", x"7F", x"00", x"C0", x"F9", x"F3", x"E1", x"FC", x"9C", x"C1", x"FF", x"3F", x"06", x"0C", x"1E", x"03", x"63", x"3E", x"00", x"F1", x"E1", x"C9", x"99", x"80", x"F9", x"F9", x"FF", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"81", x"9F", x"81", x"FC", x"FC", x"9C", x"C1", x"FF", x"7E", x"60", x"7E", x"03", x"03", x"63", x"3E", x"00", x"E1", x"CF", x"9F", x"81", x"9C", x"9C", x"C1", x"FF", x"1E", x"30", x"60", x"7E", x"63", x"63", x"3E", x"00", 
															x"80", x"9C", x"F9", x"F3", x"E7", x"E7", x"E7", x"FF", x"7F", x"63", x"06", x"0C", x"18", x"18", x"18", x"00", x"C3", x"9D", x"8D", x"C3", x"B0", x"BC", x"C1", x"FF", x"3C", x"62", x"72", x"3C", x"4F", x"43", x"3E", x"00", x"C1", x"9C", x"9C", x"C0", x"FC", x"F9", x"C3", x"FF", x"3E", x"63", x"63", x"3F", x"03", x"06", x"3C", x"00", x"FF", x"FF", x"FF", x"FF", x"E3", x"C9", x"9C", x"9C", x"00", x"00", x"00", x"00", x"1C", x"36", x"63", x"63", x"FF", x"FF", x"FF", x"FF", x"F3", x"E3", x"F3", x"F3", x"00", x"00", x"00", x"00", x"0C", x"1C", x"0C", x"0C", x"FF", x"FF", x"FF", x"FF", x"C1", x"9C", x"F8", x"E1", x"00", x"00", x"00", x"00", x"3E", x"63", x"07", x"1E", x"FF", x"FF", x"FF", x"FF", x"C0", x"F9", x"F3", x"E1", x"00", x"00", x"00", x"00", x"3F", x"06", x"0C", x"1E", x"FF", x"FF", x"FF", x"FF", x"F1", x"E1", x"C9", x"99", x"00", x"00", x"00", x"00", x"0E", x"1E", x"36", x"66", 
															x"FF", x"FF", x"FF", x"FF", x"81", x"9F", x"81", x"FC", x"00", x"00", x"00", x"00", x"7E", x"60", x"7E", x"03", x"FF", x"FF", x"FF", x"FF", x"E1", x"CF", x"9F", x"81", x"00", x"00", x"00", x"00", x"1E", x"30", x"60", x"7E", x"FF", x"FF", x"FF", x"FF", x"80", x"9C", x"F9", x"F3", x"00", x"00", x"00", x"00", x"7F", x"63", x"06", x"0C", x"FF", x"FF", x"FF", x"FF", x"C3", x"9D", x"8D", x"C3", x"00", x"00", x"00", x"00", x"3C", x"62", x"72", x"3C", x"FF", x"FF", x"FF", x"FF", x"C1", x"9C", x"9C", x"C0", x"00", x"00", x"00", x"00", x"3E", x"63", x"63", x"3F", x"9C", x"C9", x"E3", x"FF", x"FF", x"FF", x"FF", x"FF", x"63", x"36", x"1C", x"00", x"00", x"00", x"00", x"00", x"F3", x"F3", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"0C", x"0C", x"3F", x"00", x"00", x"00", x"00", x"00", x"C3", x"8F", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"3C", x"70", x"7F", x"00", x"00", x"00", x"00", x"00", 
															x"FC", x"9C", x"C1", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", x"63", x"3E", x"00", x"00", x"00", x"00", x"00", x"80", x"F9", x"F9", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"FC", x"9C", x"C1", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", x"63", x"3E", x"00", x"00", x"00", x"00", x"00", x"9C", x"9C", x"C1", x"FF", x"FF", x"FF", x"FF", x"FF", x"63", x"63", x"3E", x"00", x"00", x"00", x"00", x"00", x"E7", x"E7", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"B0", x"BC", x"C1", x"FF", x"FF", x"FF", x"FF", x"FF", x"4F", x"43", x"3E", x"00", x"00", x"00", x"00", x"00", x"FC", x"F9", x"C3", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", x"06", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"FF", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"81", x"81", x"81", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"7E", x"7E", x"7E", x"7E", x"00", x"7E", x"7E", x"7E", x"FF", x"FF", x"FF", x"FF", x"FF", x"81", x"81", x"81", x"7E", x"7E", x"7E", x"7E", x"00", x"7E", x"7E", x"7E", x"81", x"81", x"81", x"81", x"FF", x"81", x"81", x"81", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"81", x"81", x"81", x"FF", x"00", x"00", x"00", x"00", x"B9", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B9", x"46", x"49", x"49", x"49", x"49", x"49", x"49", x"46", x"99", x"66", x"E6", x"96", x"E6", x"E6", x"66", x"99", x"66", x"99", x"19", x"69", x"19", x"19", x"99", x"66", 
															x"09", x"76", x"76", x"16", x"E6", x"E6", x"E6", x"19", x"F6", x"89", x"89", x"E9", x"19", x"19", x"19", x"E6", x"FF", x"FF", x"FF", x"FF", x"B9", x"B6", x"B6", x"B6", x"00", x"00", x"00", x"00", x"46", x"49", x"49", x"49", x"B6", x"B6", x"B6", x"B9", x"FF", x"FF", x"FF", x"FF", x"49", x"49", x"49", x"46", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"99", x"66", x"E6", x"96", x"00", x"00", x"00", x"00", x"66", x"99", x"19", x"69", x"E6", x"E6", x"66", x"99", x"FF", x"FF", x"FF", x"FF", x"19", x"19", x"99", x"66", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"09", x"76", x"76", x"16", x"00", x"00", x"00", x"00", x"F6", x"89", x"89", x"E9", x"E6", x"E6", x"E6", x"19", x"FF", x"FF", x"FF", x"FF", x"19", x"19", x"19", x"E6", x"00", x"00", x"00", x"00", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"40", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", 
															x"DF", x"DF", x"DF", x"C0", x"FF", x"FF", x"FF", x"FF", x"E0", x"E0", x"E0", x"FF", x"FF", x"7F", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"02", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"FB", x"FB", x"FB", x"03", x"FF", x"FF", x"FF", x"FF", x"07", x"07", x"07", x"FF", x"FF", x"FE", x"00", x"00", x"FF", x"FF", x"F7", x"38", x"FF", x"FF", x"F7", x"F7", x"00", x"00", x"18", x"FF", x"FF", x"FF", x"18", x"18", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"18", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"38", x"44", x"82", x"80", x"8E", x"82", x"44", x"38", x"38", x"44", x"82", x"80", x"8E", x"82", x"44", x"38", x"38", x"44", x"82", x"80", x"8E", x"82", x"44", x"38", 
															x"FF", x"FF", x"FF", x"FF", x"F8", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"0F", x"08", x"08", x"08", x"08", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"00", x"F0", x"10", x"10", x"10", x"10", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"F8", x"F8", x"F8", x"FF", x"F8", x"F8", x"F8", x"F8", x"08", x"08", x"08", x"0F", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"FF", x"1F", x"1F", x"1F", x"1F", x"10", x"10", x"10", x"F0", x"10", x"10", x"10", x"10", 
															x"F8", x"F8", x"F8", x"FF", x"FF", x"FF", x"FF", x"FF", x"08", x"08", x"08", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"FF", x"FF", x"FF", x"FF", x"FF", x"10", x"10", x"10", x"F0", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"E0", x"60", x"70", x"38", x"1E", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"E0", x"07", x"07", x"0E", x"0E", x"1C", x"1C", x"38", x"F0", x"00", x"00", x"01", x"01", x"03", x"03", x"07", x"0F", x"18", x"10", x"10", x"30", x"20", x"20", x"60", x"40", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"80", x"80", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"83", x"C0", x"60", x"38", x"0F", x"01", x"F0", x"F8", x"7C", x"3F", x"1F", x"07", x"00", x"00", 
															x"01", x"FF", x"FF", x"FE", x"00", x"00", x"01", x"FF", x"00", x"00", x"00", x"01", x"FF", x"FF", x"FE", x"00", x"E0", x"C1", x"83", x"06", x"0C", x"38", x"E0", x"00", x"1F", x"3E", x"7C", x"F8", x"F0", x"C0", x"00", x"00", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"2F", x"68", x"68", x"AE", x"A1", x"F1", x"21", x"2E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"89", x"89", x"E9", x"19", x"19", x"19", x"E6", x"3C", x"20", x"20", x"38", x"04", x"04", x"04", x"38", x"3C", x"20", x"20", x"38", x"04", x"04", x"04", x"38", x"46", x"49", x"49", x"49", x"49", x"49", x"49", x"46", x"46", x"49", x"49", x"49", x"49", x"49", x"49", x"46", x"4F", x"48", x"48", x"4E", x"41", x"41", x"41", x"4E", x"4F", x"48", x"48", x"4E", x"41", x"41", x"41", x"4E", 
															x"66", x"99", x"19", x"19", x"29", x"49", x"89", x"F6", x"66", x"99", x"19", x"19", x"29", x"49", x"89", x"F6", x"6F", x"98", x"18", x"1E", x"21", x"41", x"81", x"FE", x"6F", x"98", x"18", x"1E", x"21", x"41", x"81", x"FE", x"66", x"99", x"19", x"69", x"19", x"19", x"99", x"66", x"66", x"99", x"19", x"69", x"19", x"19", x"99", x"66", x"6F", x"98", x"18", x"6E", x"11", x"11", x"91", x"6E", x"6F", x"98", x"18", x"6E", x"11", x"11", x"91", x"6E", x"26", x"69", x"69", x"A9", x"A9", x"F9", x"29", x"26", x"26", x"69", x"69", x"A9", x"A9", x"F9", x"29", x"26", x"2F", x"68", x"68", x"AE", x"A1", x"F1", x"21", x"2E", x"2F", x"68", x"68", x"AE", x"A1", x"F1", x"21", x"2E", x"F6", x"89", x"89", x"E9", x"19", x"19", x"19", x"E6", x"F6", x"89", x"89", x"E9", x"19", x"19", x"19", x"E6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
	
	constant TENNIS_CHR_ROM : CHR_ROM_ARRAY := (x"38", x"68", x"54", x"6C", x"54", x"6C", x"3C", x"0C", x"00", x"20", x"10", x"28", x"10", x"28", x"00", x"00", x"00", x"00", x"00", x"3C", x"7F", x"78", x"72", x"60", x"00", x"00", x"00", x"00", x"00", x"06", x"0C", x"1F", x"04", x"04", x"00", x"02", x"02", x"00", x"00", x"00", x"00", x"02", x"07", x"05", x"05", x"00", x"00", x"00", x"03", x"00", x"06", x"0F", x"1F", x"0F", x"07", x"07", x"00", x"03", x"07", x"0E", x"1F", x"1F", x"3D", x"FB", x"00", x"00", x"40", x"60", x"E0", x"E0", x"C0", x"80", x"F0", x"E0", x"C0", x"E0", x"60", x"F0", x"F0", x"BE", x"0F", x"1F", x"1F", x"3F", x"3F", x"3F", x"1E", x"00", x"FF", x"FF", x"47", x"00", x"00", x"00", x"00", x"1E", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"3E", x"08", x"00", x"00", x"40", x"E0", x"F0", x"70", x"00", x"00", x"00", x"00", x"20", x"70", x"78", x"3C", x"0E", x"0E", x"1E", x"1C", x"18", x"40", x"78", x"3C", 
															x"00", x"C0", x"E0", x"70", x"30", x"00", x"00", x"00", x"70", x"A0", x"C0", x"70", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7F", x"78", x"72", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"0C", x"06", x"06", x"00", x"0C", x"1E", x"3F", x"3F", x"0F", x"01", x"01", x"07", x"0F", x"1D", x"3E", x"3F", x"3B", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"80", x"F0", x"E0", x"C0", x"00", x"C0", x"E0", x"F0", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"1B", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"07", x"0F", x"0F", x"1F", x"3F", x"BF", x"BE", x"3C", x"3F", x"7F", x"7F", x"FE", x"C0", x"40", x"41", x"00", x"36", x"6A", x"56", x"6A", x"54", x"2C", x"18", x"00", x"10", x"28", x"14", x"28", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"E0", x"F0", x"78", x"1C", x"1C", x"3C", x"38", x"30", x"80", x"F0", x"78", 
															x"00", x"00", x"3C", x"3E", x"30", x"00", x"00", x"00", x"30", x"30", x"0C", x"3E", x"30", x"00", x"00", x"00", x"0C", x"00", x"18", x"1E", x"3E", x"3E", x"3F", x"7C", x"03", x"0F", x"16", x"18", x"3D", x"3F", x"3F", x"6F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"80", x"00", x"00", x"00", x"C0", x"80", x"00", x"1E", x"1E", x"1F", x"3F", x"3F", x"3F", x"39", x"00", x"1D", x"1F", x"07", x"00", x"00", x"00", x"06", x"1E", x"00", x"00", x"00", x"00", x"86", x"83", x"00", x"00", x"C0", x"E0", x"F0", x"7C", x"18", x"6C", x"F0", x"F0", x"78", x"AC", x"D6", x"AA", x"56", x"6C", x"18", x"00", x"00", x"28", x"54", x"28", x"14", x"08", x"00", x"00", x"00", x"00", x"00", x"60", x"F0", x"E0", x"70", x"78", x"0E", x"0E", x"1E", x"5C", x"E8", x"E0", x"70", x"78", x"00", x"3C", x"38", x"30", x"00", x"00", x"00", x"00", x"30", x"0C", x"38", x"30", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"3E", x"7F", x"7C", x"7C", x"7C", x"00", x"00", x"00", x"00", x"00", x"02", x"02", x"02", x"30", x"58", x"AC", x"D4", x"AC", x"D4", x"E8", x"30", x"00", x"10", x"28", x"50", x"28", x"50", x"20", x"00", x"0F", x"00", x"0F", x"3F", x"7F", x"7F", x"3F", x"3F", x"00", x"07", x"0F", x"3F", x"7F", x"7F", x"7F", x"7F", x"00", x"01", x"03", x"C0", x"C0", x"C0", x"80", x"00", x"C0", x"80", x"04", x"FE", x"FE", x"F0", x"80", x"00", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"0E", x"00", x"0F", x"0F", x"01", x"00", x"00", x"00", x"01", x"0F", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"C0", x"80", x"80", x"00", x"40", x"60", x"70", x"70", x"00", x"00", x"00", x"78", x"78", x"70", x"38", x"38", x"07", x"07", x"0F", x"66", x"74", x"70", x"38", x"38", x"70", x"D0", x"A8", x"D9", x"AB", x"DB", x"7F", x"07", x"00", x"40", x"20", x"50", x"20", x"50", x"00", x"00", 
															x"00", x"00", x"00", x"E0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"01", x"01", x"0F", x"1F", x"3F", x"0F", x"0F", x"07", x"00", x"01", x"0F", x"1F", x"3F", x"7F", x"7F", x"3F", x"E0", x"B0", x"F0", x"F0", x"F0", x"E0", x"E0", x"C0", x"10", x"F8", x"FC", x"F8", x"F0", x"E0", x"E0", x"C0", x"0F", x"0F", x"1F", x"1F", x"1F", x"0F", x"04", x"00", x"0F", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"C0", x"C0", x"80", x"80", x"80", x"80", x"80", x"00", x"C0", x"C0", x"00", x"40", x"60", x"60", x"70", x"70", x"00", x"00", x"02", x"06", x"0F", x"0D", x"08", x"00", x"0F", x"07", x"03", x"07", x"0E", x"0F", x"0F", x"07", x"D8", x"30", x"60", x"61", x"F9", x"F1", x"F3", x"74", x"18", x"FE", x"BF", x"BE", x"7E", x"F2", x"F0", x"F3", x"60", x"D0", x"A8", x"58", x"A8", x"58", x"B0", x"60", x"00", x"40", x"20", x"50", x"A0", x"50", x"20", x"00", 
															x"00", x"00", x"01", x"03", x"03", x"01", x"01", x"00", x"03", x"01", x"00", x"00", x"04", x"0E", x"1E", x"1C", x"04", x"20", x"C8", x"FC", x"FC", x"FC", x"78", x"00", x"FA", x"D8", x"30", x"00", x"00", x"00", x"00", x"78", x"00", x"00", x"00", x"03", x"07", x"07", x"01", x"00", x"0F", x"07", x"03", x"03", x"07", x"07", x"07", x"07", x"60", x"60", x"18", x"3C", x"78", x"F0", x"F0", x"F0", x"80", x"80", x"F8", x"FC", x"BE", x"7E", x"FE", x"FE", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"07", x"03", x"00", x"00", x"02", x"07", x"0F", x"0F", x"78", x"18", x"10", x"31", x"C3", x"FD", x"7D", x"79", x"FE", x"FE", x"FE", x"CC", x"3C", x"00", x"80", x"00", x"00", x"E0", x"50", x"A8", x"58", x"A8", x"D8", x"70", x"00", x"00", x"40", x"A0", x"50", x"A0", x"50", x"00", x"0C", x"00", x"06", x"2F", x"7F", x"3F", x"27", x"23", x"F0", x"7C", x"1E", x"37", x"6F", x"7F", x"FF", x"FF", 
															x"00", x"0F", x"1A", x"35", x"2A", x"35", x"1B", x"0E", x"00", x"00", x"0A", x"15", x"0A", x"14", x"0A", x"00", x"00", x"00", x"00", x"21", x"E1", x"81", x"80", x"00", x"0B", x"0F", x"3F", x"1C", x"1A", x"06", x"07", x"0E", x"30", x"70", x"F8", x"F8", x"F8", x"F8", x"B8", x"00", x"F0", x"F0", x"E0", x"00", x"00", x"00", x"40", x"78", x"70", x"68", x"D4", x"AC", x"D4", x"AC", x"54", x"3C", x"00", x"20", x"50", x"28", x"50", x"28", x"10", x"00", x"60", x"20", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"18", x"1F", x"1D", x"0F", x"07", x"03", x"00", x"3C", x"00", x"7C", x"FE", x"FE", x"FE", x"FE", x"3E", x"C0", x"78", x"FC", x"FE", x"FE", x"FE", x"FE", x"3E", x"0E", x"1B", x"15", x"9B", x"D5", x"FE", x"C0", x"C0", x"00", x"0A", x"04", x"0A", x"04", x"00", x"00", x"30", x"80", x"C0", x"E0", x"F0", x"E0", x"E0", x"E0", x"E0", x"70", x"E0", x"F0", x"F8", x"F8", x"F8", x"E0", x"E0", 
															x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F8", x"E2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"03", x"03", x"03", x"07", x"0F", x"0F", x"1F", x"1F", x"00", x"00", x"00", x"07", x"0F", x"0F", x"1F", x"1F", x"E7", x"C5", x"C7", x"E5", x"F3", x"FE", x"FC", x"F8", x"12", x"30", x"32", x"E0", x"FE", x"F8", x"F8", x"FC", x"1F", x"1F", x"1F", x"3F", x"3F", x"3F", x"3F", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"00", x"00", x"00", x"F0", x"C0", x"80", x"80", x"80", x"C0", x"C0", x"80", x"DC", x"FC", x"98", x"80", x"00", x"00", x"20", x"60", x"01", x"00", x"00", x"00", x"00", x"30", x"70", x"78", x"1C", x"1C", x"3C", x"38", x"38", x"00", x"70", x"78", x"00", x"00", x"00", x"00", x"00", x"60", x"70", x"78", x"F0", x"F0", x"F0", x"70", x"60", x"00", x"70", x"78", 
															x"00", x"00", x"00", x"00", x"00", x"7C", x"FE", x"F9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"1F", x"1E", x"1E", x"3F", x"7F", x"7F", x"7F", x"FF", x"00", x"01", x"01", x"3F", x"7F", x"7F", x"7F", x"FF", x"70", x"50", x"70", x"50", x"90", x"F0", x"E0", x"C0", x"A0", x"80", x"A0", x"00", x"E0", x"C0", x"C0", x"E0", x"3F", x"3F", x"3F", x"3F", x"7F", x"7F", x"7F", x"3F", x"3F", x"3F", x"3F", x"01", x"00", x"00", x"00", x"00", x"E0", x"80", x"00", x"00", x"80", x"C0", x"C0", x"80", x"B8", x"F8", x"30", x"00", x"00", x"00", x"00", x"40", x"02", x"00", x"00", x"00", x"00", x"60", x"70", x"78", x"39", x"39", x"38", x"70", x"70", x"00", x"70", x"78", x"00", x"00", x"00", x"00", x"00", x"60", x"70", x"78", x"E0", x"E0", x"E0", x"60", x"60", x"00", x"70", x"78", x"00", x"01", x"01", x"01", x"00", x"1C", x"1E", x"0F", x"1F", x"0E", x"07", x"0F", x"0E", x"10", x"1E", x"0F", 
															x"00", x"00", x"80", x"C0", x"C0", x"00", x"00", x"00", x"C0", x"C0", x"00", x"C0", x"C0", x"00", x"00", x"00", x"02", x"02", x"C0", x"E0", x"60", x"60", x"20", x"00", x"0D", x"1D", x"BE", x"D8", x"60", x"60", x"20", x"00", x"0F", x"1F", x"1F", x"3F", x"3F", x"3F", x"1E", x"01", x"FF", x"FF", x"43", x"00", x"00", x"00", x"01", x"1E", x"80", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"9F", x"0C", x"00", x"00", x"00", x"00", x"80", x"C0", x"0F", x"1F", x"1F", x"1F", x"1F", x"1F", x"0F", x"04", x"FF", x"FF", x"47", x"00", x"00", x"00", x"00", x"0B", x"80", x"00", x"00", x"80", x"80", x"C0", x"00", x"00", x"9F", x"04", x"00", x"00", x"00", x"00", x"C0", x"C0", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"03", x"01", x"00", x"00", x"00", x"00", x"01", x"03", x"04", x"20", x"CC", x"FC", x"FC", x"FC", x"78", x"80", x"FA", x"D8", x"F8", x"00", x"00", x"00", x"80", x"78", 
															x"00", x"00", x"00", x"01", x"01", x"03", x"00", x"00", x"03", x"01", x"00", x"00", x"00", x"00", x"03", x"03", x"04", x"20", x"C8", x"F8", x"F8", x"F8", x"F0", x"20", x"FA", x"D8", x"F0", x"00", x"00", x"00", x"00", x"D0", x"00", x"00", x"3C", x"7F", x"78", x"72", x"60", x"60", x"00", x"00", x"00", x"00", x"06", x"0C", x"1F", x"1E", x"00", x"0E", x"1F", x"3F", x"0F", x"0F", x"07", x"07", x"03", x"0F", x"1E", x"3F", x"3F", x"7F", x"77", x"67", x"00", x"78", x"78", x"F8", x"E0", x"E0", x"E0", x"C0", x"C0", x"FF", x"FF", x"7F", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"23", x"23", x"23", x"20", x"70", x"39", x"71", x"70", x"50", x"00", x"00", x"03", x"03", x"F0", x"F0", x"F8", x"FC", x"F8", x"E0", x"00", x"00", x"F0", x"C0", x"00", x"00", x"04", x"1E", x"DE", x"CE", 
															x"D8", x"A8", x"D8", x"A8", x"DB", x"77", x"07", x"07", x"53", x"23", x"53", x"23", x"50", x"07", x"07", x"07", x"00", x"0C", x"0E", x"0F", x"00", x"00", x"80", x"80", x"8C", x"80", x"0E", x"0F", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"03", x"07", x"0E", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"C0", x"80", x"00", x"40", x"00", x"01", x"0B", x"0E", x"06", x"06", x"C6", x"AE", x"EE", x"00", x"02", x"00", x"00", x"0C", x"08", x"08", x"38", x"00", x"04", x"0F", x"0F", x"03", x"01", x"01", x"00", x"0E", x"0E", x"07", x"0E", x"3F", x"1F", x"1F", x"1F", x"01", x"01", x"00", x"0D", x"BE", x"FF", x"FF", x"FF", x"00", x"10", x"38", x"38", x"38", x"F0", x"F0", x"E0", x"EE", x"FC", x"FC", x"F8", x"F8", x"30", x"F0", x"E0", x"58", x"A8", x"D8", x"A8", x"D8", x"B0", x"70", x"00", x"10", x"20", x"50", x"20", x"50", x"20", x"00", x"00", 
															x"07", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"1F", x"07", x"0F", x"0F", x"0F", x"03", x"00", x"00", x"00", x"E0", x"C0", x"C0", x"C0", x"E0", x"E0", x"C0", x"80", x"E0", x"C0", x"C0", x"80", x"80", x"10", x"38", x"78", x"0E", x"00", x"00", x"00", x"00", x"18", x"1C", x"3E", x"01", x"0F", x"07", x"07", x"0F", x"06", x"18", x"3E", x"00", x"00", x"38", x"3C", x"00", x"00", x"00", x"00", x"38", x"30", x"88", x"BC", x"00", x"00", x"00", x"00", x"1E", x"2B", x"35", x"2A", x"35", x"0E", x"00", x"00", x"00", x"0A", x"15", x"0A", x"04", x"00", x"00", x"00", x"00", x"00", x"E0", x"80", x"00", x"00", x"00", x"00", x"00", x"1C", x"1E", x"1F", x"07", x"03", x"01", x"01", x"00", x"00", x"30", x"60", x"40", x"28", x"20", x"60", x"00", x"00", x"00", x"00", x"B8", x"D4", x"FC", x"FC", x"F8", x"F8", x"7C", x"7C", x"7C", x"7C", x"7C", x"FC", x"FE", x"FC", x"7C", x"7E", x"7F", x"7E", x"7C", x"FC", 
															x"1F", x"3F", x"7F", x"7E", x"7E", x"0E", x"04", x"00", x"1F", x"07", x"01", x"00", x"00", x"31", x"7B", x"7B", x"00", x"00", x"00", x"18", x"1C", x"38", x"1C", x"0E", x"07", x"0F", x"0E", x"06", x"10", x"38", x"1C", x"0E", x"00", x"00", x"70", x"78", x"00", x"00", x"00", x"00", x"60", x"60", x"10", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"58", x"AC", x"D4", x"00", x"00", x"00", x"00", x"00", x"10", x"28", x"50", x"AC", x"D4", x"68", x"30", x"10", x"10", x"10", x"00", x"28", x"50", x"20", x"00", x"00", x"00", x"00", x"38", x"00", x"00", x"1E", x"3F", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"00", x"00", x"01", x"07", x"1F", x"7F", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"80", x"38", x"30", x"70", x"F0", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"01", x"03", x"03", x"00", x"00", x"00", x"00", 
															x"FF", x"7F", x"FE", x"FC", x"FC", x"F8", x"F8", x"F8", x"FF", x"FF", x"FE", x"FC", x"FC", x"F8", x"08", x"00", x"01", x"01", x"00", x"06", x"0E", x"1E", x"1E", x"18", x"00", x"00", x"00", x"06", x"0E", x"1D", x"1D", x"18", x"F8", x"F8", x"88", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"70", x"F0", x"F0", x"E0", x"E0", x"C0", x"60", x"60", x"70", x"38", x"00", x"00", x"00", x"00", x"00", x"60", x"70", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"1F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"3F", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"3F", x"1F", x"3F", x"3F", x"3F", x"3F", x"3E", x"7F", x"3F", x"7F", x"FF", x"FF", x"3F", x"3F", x"00", x"00", x"F0", x"C0", x"80", x"82", x"1E", x"2B", x"35", x"1E", x"FE", x"C7", x"87", x"80", x"00", x"0A", x"14", x"00", 
															x"7F", x"7F", x"30", x"00", x"40", x"E0", x"E0", x"E0", x"00", x"00", x"0F", x"37", x"57", x"DF", x"DE", x"DC", x"D8", x"D8", x"1C", x"0E", x"00", x"00", x"00", x"00", x"C0", x"D8", x"1C", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"03", x"07", x"07", x"07", x"7F", x"DF", x"01", x"07", x"0F", x"1F", x"1F", x"07", x"00", x"50", x"F8", x"F8", x"FC", x"FC", x"F8", x"E0", x"C0", x"E0", x"F4", x"F8", x"FC", x"FC", x"FC", x"FC", x"30", x"00", x"1A", x"15", x"1B", x"0E", x"00", x"00", x"00", x"00", x"0A", x"05", x"0A", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"E1", x"00", x"00", x"70", x"78", x"78", x"01", x"01", x"1F", x"EF", x"6F", x"6F", x"E6", x"F0", x"70", x"F0", x"E0", x"F0", x"00", x"00", x"00", x"00", x"F0", x"30", x"C0", x"F0", x"00", x"00", x"00", x"00", 
															x"03", x"00", x"39", x"7B", x"1F", x"0F", x"1F", x"0F", x"3C", x"1F", x"3E", x"7D", x"7B", x"FE", x"FE", x"7C", x"70", x"E0", x"E0", x"D0", x"B0", x"50", x"B0", x"50", x"70", x"FC", x"9E", x"4E", x"27", x"47", x"A5", x"41", x"01", x"00", x"01", x"03", x"03", x"01", x"00", x"00", x"1E", x"0E", x"00", x"00", x"04", x"06", x"0F", x"0E", x"F8", x"F8", x"F8", x"FC", x"FC", x"FC", x"BC", x"00", x"40", x"F8", x"E0", x"00", x"00", x"00", x"00", x"38", x"18", x"2C", x"57", x"6C", x"54", x"6C", x"58", x"30", x"01", x"09", x"10", x"28", x"10", x"28", x"10", x"00", x"00", x"00", x"06", x"0E", x"0F", x"03", x"03", x"03", x"EF", x"F7", x"BF", x"1F", x"0E", x"03", x"03", x"03", x"C0", x"3C", x"70", x"F0", x"F8", x"F0", x"F0", x"F0", x"00", x"FC", x"BE", x"7F", x"FF", x"F3", x"F7", x"F3", x"01", x"01", x"01", x"03", x"01", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"06", x"06", x"0F", x"0E", 
															x"F0", x"F8", x"F8", x"F8", x"F8", x"F8", x"78", x"00", x"F0", x"F8", x"E0", x"00", x"00", x"00", x"00", x"70", x"80", x"C0", x"40", x"0F", x"1F", x"07", x"07", x"07", x"00", x"30", x"38", x"70", x"00", x"08", x"08", x"08", x"00", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"3C", x"22", x"60", x"70", x"40", x"01", x"0F", x"D8", x"7C", x"3E", x"7E", x"7F", x"7F", x"FF", x"7F", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"C0", x"E0", x"E0", x"E0", x"C0", x"00", x"E0", x"F0", x"00", x"1C", x"34", x"2A", x"36", x"2A", x"36", x"1C", x"00", x"00", x"10", x"08", x"14", x"08", x"14", x"00", x"04", x"06", x"02", x"E0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"03", x"03", x"07", x"06", x"0E", x"E0", x"B0", x"F8", x"F8", x"F0", x"E0", x"E0", x"C0", x"0E", x"FC", x"FC", x"F8", x"F0", x"E0", x"E0", x"C0", 
															x"00", x"00", x"00", x"0C", x"0A", x"16", x"1A", x"14", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"00", x"1C", x"11", x"17", x"00", x"02", x"00", x"02", x"03", x"00", x"00", x"00", x"1B", x"19", x"0B", x"0F", x"0F", x"00", x"C0", x"E0", x"20", x"A0", x"00", x"00", x"70", x"00", x"00", x"00", x"C0", x"40", x"E0", x"E0", x"F0", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"01", x"00", x"0F", x"0F", x"0C", x"00", x"01", x"F8", x"B8", x"18", x"18", x"38", x"7C", x"FC", x"4C", x"F8", x"F8", x"E8", x"F8", x"F8", x"30", x"00", x"B0", x"00", x"00", x"00", x"03", x"07", x"00", x"00", x"00", x"03", x"03", x"03", x"00", x"07", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"0C", x"0C", x"18", x"00", x"B8", x"70", x"70", x"38", x"34", x"0C", x"18", x"00", x"00", x"00", x"1C", x"7E", x"02", x"2A", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"14", x"3E", x"1E", 
															x"00", x"70", x"A8", x"D8", x"A0", x"70", x"00", x"00", x"00", x"00", x"20", x"50", x"20", x"00", x"00", x"00", x"81", x"C1", x"61", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"17", x"3F", x"3C", x"01", x"01", x"00", x"30", x"78", x"C8", x"C8", x"08", x"0C", x"7C", x"7C", x"F0", x"F8", x"F8", x"F8", x"F8", x"FC", x"78", x"80", x"00", x"00", x"00", x"03", x"07", x"00", x"00", x"00", x"01", x"01", x"03", x"00", x"07", x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"C0", x"B8", x"B8", x"30", x"38", x"18", x"04", x"3C", x"00", x"00", x"38", x"FC", x"04", x"54", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"28", x"7C", x"3C", x"00", x"00", x"30", x"50", x"6C", x"54", x"38", x"00", x"00", x"00", x"00", x"10", x"28", x"10", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"B0", x"60", x"01", x"01", x"01", x"01", x"03", x"0F", x"0E", x"00", 
															x"9E", x"F8", x"F0", x"7C", x"78", x"70", x"78", x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"7E", x"06", x"00", x"0C", x"00", x"00", x"E0", x"E0", x"00", x"06", x"0F", x"33", x"77", x"67", x"86", x"E6", x"06", x"00", x"0F", x"00", x"78", x"F8", x"88", x"50", x"00", x"01", x"F9", x"00", x"00", x"00", x"70", x"A8", x"F8", x"70", x"FA", x"30", x"58", x"A8", x"D8", x"B0", x"E0", x"80", x"00", x"00", x"10", x"20", x"50", x"20", x"00", x"00", x"00", x"C0", x"C4", x"44", x"7C", x"78", x"F8", x"FC", x"FC", x"FF", x"FE", x"7C", x"7E", x"7F", x"7A", x"00", x"00", x"18", x"00", x"40", x"40", x"60", x"00", x"0E", x"07", x"27", x"37", x"73", x"77", x"66", x"06", x"08", x"07", x"00", x"03", x"37", x"5C", x"6D", x"50", x"38", x"07", x"00", x"00", x"00", x"13", x"2A", x"17", x"07", x"07", x"00", x"80", x"E0", x"00", x"40", x"00", x"00", x"80", x"00", x"00", x"00", x"C0", x"80", x"C0", x"80", x"C0", 
															x"0F", x"1F", x"1F", x"1E", x"3E", x"3E", x"3E", x"36", x"0F", x"1F", x"1F", x"1E", x"1E", x"0C", x"01", x"09", x"C0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"03", x"07", x"04", x"05", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"02", x"07", x"07", x"00", x"00", x"80", x"E6", x"0D", x"4B", x"0D", x"0B", x"00", x"00", x"00", x"00", x"C4", x"82", x"C4", x"82", x"0F", x"1F", x"1C", x"1C", x"1E", x"3E", x"3E", x"3E", x"0F", x"1F", x"1F", x"1B", x"1F", x"3E", x"1E", x"01", x"0E", x"88", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"80", x"98", x"E8", x"F0", x"30", x"00", x"00", x"00", x"00", x"1C", x"3F", x"20", x"2A", x"00", x"60", x"00", x"00", x"00", x"00", x"1E", x"14", x"3E", x"7C", x"F4", x"DE", x"8C", x"0C", x"44", x"E0", x"F2", x"FC", x"FC", x"FE", x"FE", x"7E", x"7E", x"FE", x"0D", x"03", 
															x"00", x"00", x"38", x"D4", x"6C", x"54", x"38", x"00", x"00", x"00", x"00", x"10", x"28", x"10", x"00", x"00", x"00", x"00", x"18", x"34", x"2C", x"34", x"2C", x"18", x"00", x"00", x"00", x"10", x"08", x"10", x"08", x"00", x"08", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"0C", x"0F", x"0F", x"0D", x"07", x"03", x"00", x"00", x"38", x"7C", x"44", x"28", x"00", x"00", x"18", x"00", x"00", x"00", x"38", x"54", x"7C", x"38", x"F8", x"1C", x"9C", x"FC", x"F8", x"F8", x"7C", x"FC", x"FC", x"FC", x"FC", x"EC", x"F8", x"F8", x"78", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"02", x"15", x"03", x"00", x"00", x"00", x"00", x"00", x"3C", x"2A", x"3C", x"06", x"0F", x"03", x"03", x"01", x"00", x"00", x"03", x"07", x"0F", x"0F", x"0F", x"0F", x"07", x"03", x"00", x"38", x"F8", x"F8", x"60", x"80", x"80", x"58", x"F8", x"C8", x"98", x"98", x"B8", x"78", x"70", x"F0", x"E0", 
															x"07", x"01", x"00", x"00", x"00", x"00", x"06", x"0E", x"00", x"06", x"07", x"0E", x"0E", x"06", x"00", x"0E", x"F8", x"48", x"00", x"00", x"00", x"00", x"60", x"70", x"00", x"30", x"70", x"30", x"30", x"70", x"00", x"70", x"0C", x"1F", x"07", x"06", x"03", x"01", x"08", x"0F", x"0F", x"1F", x"1F", x"1F", x"1E", x"0E", x"0F", x"03", x"70", x"F0", x"F0", x"C0", x"00", x"00", x"80", x"E0", x"90", x"30", x"30", x"70", x"F0", x"E0", x"C0", x"80", x"1F", x"12", x"00", x"00", x"00", x"00", x"06", x"0E", x"00", x"0C", x"0E", x"0C", x"0C", x"06", x"00", x"0E", x"E0", x"80", x"00", x"00", x"00", x"00", x"60", x"70", x"00", x"60", x"E0", x"F0", x"70", x"60", x"00", x"70", x"00", x"00", x"01", x"01", x"03", x"00", x"00", x"00", x"01", x"01", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"B0", x"30", x"60", x"00", x"00", x"E0", x"C0", x"E0", x"D0", x"30", x"60", x"00", x"00", 
															x"00", x"00", x"00", x"07", x"07", x"00", x"00", x"00", x"01", x"01", x"01", x"06", x"07", x"00", x"00", x"00", x"00", x"04", x"0C", x"8C", x"98", x"80", x"00", x"00", x"D0", x"BC", x"B4", x"0C", x"98", x"80", x"00", x"00", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"01", x"06", x"07", x"07", x"00", x"00", x"00", x"F8", x"B8", x"18", x"18", x"3C", x"7C", x"9C", x"08", x"F8", x"F8", x"E8", x"F8", x"F0", x"00", x"60", x"F0", x"F8", x"B8", x"18", x"18", x"38", x"7C", x"1C", x"18", x"F8", x"F8", x"E8", x"F8", x"F0", x"00", x"E0", x"E0", x"0F", x"1F", x"1F", x"1E", x"3E", x"3E", x"38", x"10", x"0F", x"1F", x"1F", x"1E", x"0E", x"00", x"06", x"0F", x"C0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"1F", x"1E", x"1E", x"1F", x"18", x"08", x"0F", x"0F", x"1F", x"1E", x"0E", x"00", x"07", x"07", 
															x"1C", x"7E", x"02", x"2A", x"00", x"00", x"1E", x"3E", x"00", x"00", x"3C", x"14", x"3E", x"3C", x"1E", x"3E", x"00", x"00", x"01", x"03", x"35", x"5D", x"69", x"59", x"73", x"3F", x"0F", x"01", x"03", x"10", x"22", x"12", x"E0", x"60", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"E0", x"E0", x"F0", x"00", x"00", x"00", x"30", x"00", x"00", x"06", x"0E", x"00", x"00", x"00", x"07", x"06", x"06", x"00", x"0E", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"00", x"00", x"60", x"E0", x"20", x"E0", x"E0", x"E0", x"60", x"60", x"00", x"E0", x"00", x"00", x"01", x"00", x"00", x"00", x"01", x"01", x"60", x"38", x"10", x"1B", x"1B", x"1D", x"1F", x"0F", x"80", x"60", x"30", x"50", x"10", x"30", x"00", x"D0", x"00", x"80", x"C0", x"A0", x"E0", x"C0", x"E0", x"C8", x"3E", x"3E", x"3E", x"1E", x"1E", x"1F", x"3F", x"3F", x"7F", x"3F", x"3F", x"1F", x"1E", x"1F", x"1C", x"40", 
															x"00", x"40", x"7C", x"2A", x"36", x"2A", x"1C", x"00", x"C0", x"80", x"00", x"08", x"14", x"08", x"00", x"00", x"1F", x"0E", x"00", x"60", x"E0", x"00", x"06", x"1E", x"E0", x"E0", x"CE", x"0E", x"EC", x"06", x"00", x"1E", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"00", x"00", x"00", x"E0", x"50", x"B0", x"50", x"E0", x"00", x"00", x"00", x"00", x"40", x"A0", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"04", x"0F", x"0F", x"60", x"30", x"88", x"28", x"08", x"10", x"C0", x"E0", x"1C", x"C8", x"70", x"D0", x"F0", x"E0", x"E0", x"E0", x"0E", x"42", x"60", x"F0", x"F8", x"FC", x"FC", x"FC", x"7E", x"7E", x"7E", x"FC", x"F8", x"70", x"00", x"00", x"38", x"00", x"00", x"40", x"C0", x"88", x"1C", x"38", x"C4", x"DC", x"D8", x"98", x"D8", x"90", x"0C", x"38", 
															x"00", x"00", x"60", x"B0", x"D0", x"B0", x"D0", x"60", x"00", x"00", x"00", x"20", x"40", x"20", x"40", x"00", x"20", x"20", x"00", x"00", x"00", x"00", x"02", x"03", x"00", x"00", x"60", x"60", x"60", x"30", x"30", x"30", x"00", x"00", x"03", x"03", x"03", x"03", x"03", x"07", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"07", x"18", x"C4", x"94", x"C4", x"C8", x"E0", x"F0", x"38", x"60", x"B8", x"E8", x"F8", x"F0", x"F0", x"F0", x"F8", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"03", x"00", x"07", x"07", x"0F", x"07", x"00", x"00", x"0C", x"0D", x"08", x"80", x"C0", x"C0", x"C0", x"E0", x"00", x"00", x"F8", x"F8", x"D8", x"80", x"00", x"00", x"C0", x"C0", x"00", x"80", x"C0", x"C0", x"40", x"0E", x"06", x"03", x"6E", x"EE", x"A6", x"C6", x"46", x"08", x"06", x"03", x"00", x"1C", x"3F", x"21", x"28", x"02", x"E0", x"F8", x"00", x"00", x"00", x"1E", x"16", x"3C", x"FE", x"FC", 
															x"03", x"03", x"03", x"07", x"07", x"0F", x"0F", x"0F", x"03", x"03", x"03", x"07", x"07", x"03", x"00", x"00", x"C0", x"80", x"C0", x"E0", x"C0", x"C0", x"80", x"C6", x"F0", x"F8", x"F8", x"F8", x"D8", x"CC", x"8C", x"00", x"4C", x"00", x"00", x"C0", x"C0", x"C0", x"06", x"07", x"32", x"3B", x"3B", x"B7", x"B6", x"C6", x"00", x"07", x"1E", x"0D", x"0B", x"0D", x"06", x"00", x"00", x"00", x"00", x"04", x"02", x"04", x"00", x"00", x"00", x"00", x"18", x"00", x"00", x"06", x"06", x"60", x"60", x"E0", x"E4", x"EC", x"6C", x"6A", x"66", x"00", x"60", x"E0", x"00", x"06", x"8B", x"ED", x"0B", x"4D", x"0E", x"18", x"00", x"00", x"02", x"04", x"C2", x"84", x"C0", x"80", x"0F", x"1E", x"1C", x"1C", x"1F", x"3E", x"3E", x"3E", x"0F", x"1F", x"1F", x"1F", x"1F", x"1E", x"0E", x"01", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"C0", x"E0", x"00", x"00", x"80", x"80", x"C0", x"C0", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"1C", x"14", x"1C", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"08", x"14", x"1C", x"0C", x"04", x"04", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"02", x"07", x"07", x"03", x"00", x"0E", x"1F", x"11", x"0A", x"00", x"00", x"33", x"00", x"00", x"00", x"0E", x"15", x"1F", x"CE", x"FF", x"3F", x"7F", x"3F", x"3E", x"3E", x"1F", x"3F", x"3F", x"FF", x"7F", x"3F", x"3E", x"3E", x"1E", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"60", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"7C", x"7C", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"FE", x"FE", x"FE", x"FE", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"18", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"7C", x"38", x"00", x"00", x"00", x"00", x"18", x"2C", x"54", x"6C", x"54", x"6C", x"00", x"00", x"00", x"08", x"10", x"28", x"10", x"28", x"38", x"30", x"60", x"47", x"4F", x"0F", x"0F", x"0F", x"10", x"00", x"00", x"00", x"80", x"C0", x"F0", x"D0", x"07", x"0D", x"0F", x"1F", x"0F", x"07", x"07", x"03", x"78", x"7F", x"3F", x"1F", x"0F", x"07", x"07", x"03", x"80", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"10", x"38", x"6C", x"C6", x"82", x"82", x"82", x"00", x"00", x"00", x"10", x"38", x"7C", x"7C", x"7C", x"92", x"54", x"38", x"FE", x"38", x"54", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C7", x"B3", x"39", x"39", x"39", x"9B", x"C7", x"FF", x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"E7", x"C7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"83", x"39", x"F1", x"C3", x"87", x"1F", x"01", x"FF", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"81", x"F3", x"E7", x"C3", x"F9", x"39", x"83", x"FF", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"E3", x"C3", x"93", x"33", x"01", x"F3", x"F3", x"FF", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"03", x"3F", x"03", x"F9", x"F9", x"39", x"83", x"FF", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"E1", x"CF", x"9F", x"81", x"9C", x"9C", x"C1", x"FF", x"1E", x"30", x"60", x"7E", x"63", x"63", x"3E", x"00", x"01", x"39", x"F3", x"E7", x"CF", x"CF", x"CF", x"FF", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", 
															x"87", x"3B", x"1B", x"87", x"79", x"79", x"83", x"FF", x"78", x"C4", x"E4", x"78", x"86", x"86", x"7C", x"00", x"83", x"39", x"39", x"81", x"F9", x"F3", x"87", x"FF", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"C7", x"93", x"39", x"39", x"01", x"39", x"39", x"FF", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"03", x"39", x"39", x"03", x"39", x"39", x"03", x"FF", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"C3", x"99", x"3F", x"3F", x"3F", x"99", x"C3", x"FF", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"07", x"33", x"39", x"39", x"39", x"33", x"07", x"FF", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"01", x"3F", x"3F", x"03", x"3F", x"3F", x"01", x"FF", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"33", x"33", x"94", x"85", x"CD", x"CC", x"CC", x"FF", x"CC", x"CC", x"6B", x"7A", x"32", x"33", x"33", x"00", 
															x"C1", x"9F", x"3F", x"31", x"39", x"99", x"C1", x"FF", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"FF", x"FF", x"57", x"57", x"57", x"47", x"47", x"FF", x"00", x"00", x"A8", x"A8", x"A8", x"B8", x"B8", x"00", x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"20", x"00", x"00", x"00", x"00", x"8F", x"0F", x"38", x"3A", x"3A", x"08", x"88", x"FF", x"70", x"F0", x"C7", x"C5", x"C5", x"F7", x"77", x"00", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"81", x"FF", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"39", x"11", x"01", x"01", x"29", x"39", x"39", x"FF", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"39", x"19", x"09", x"01", x"21", x"31", x"39", x"FF", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", 
															x"83", x"39", x"39", x"39", x"39", x"39", x"83", x"FF", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"03", x"39", x"39", x"39", x"03", x"3F", x"3F", x"FF", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"03", x"39", x"39", x"31", x"07", x"23", x"31", x"FF", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"87", x"33", x"3F", x"83", x"F9", x"39", x"83", x"FF", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"39", x"39", x"39", x"39", x"39", x"39", x"83", x"FF", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"39", x"39", x"39", x"11", x"83", x"C7", x"EF", x"FF", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", 
															x"39", x"39", x"29", x"01", x"01", x"11", x"39", x"FF", x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"39", x"11", x"83", x"C7", x"83", x"11", x"39", x"FF", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"99", x"99", x"99", x"C3", x"E7", x"E7", x"E7", x"FF", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"FF", x"FF", x"FF", x"FF", x"9F", x"9F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"F3", x"F3", x"F3", x"F7", x"FF", x"E7", x"E7", x"FF", x"0C", x"0C", x"0C", x"08", x"00", x"18", x"18", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"93", x"93", x"F7", x"FF", x"00", x"00", x"00", x"00", x"6C", x"6C", x"08", x"00", x"FF", x"C3", x"E7", x"E7", x"E7", x"E7", x"C3", x"FF", x"00", x"3C", x"18", x"18", x"18", x"18", x"3C", x"00", x"FF", x"83", x"D7", x"D7", x"D7", x"D7", x"83", x"FF", x"00", x"7C", x"28", x"28", x"28", x"28", x"7C", x"00", x"FF", x"01", x"AB", x"AB", x"AB", x"AB", x"01", x"FF", x"00", x"FE", x"54", x"54", x"54", x"54", x"FE", x"00", x"D7", x"81", x"55", x"07", x"D3", x"55", x"01", x"D7", x"28", x"7E", x"AA", x"F8", x"2C", x"AA", x"FE", x"28", x"FF", x"FD", x"F9", x"FD", x"CF", x"CF", x"DF", x"FF", x"06", x"0F", x"0E", x"72", x"78", x"73", x"2F", x"3F", x"FF", x"FF", x"FF", x"F3", x"E5", x"F3", x"FF", x"FF", x"00", x"00", x"0C", x"1E", x"1E", x"3E", x"1E", x"00", x"FF", x"DF", x"8F", x"9F", x"F9", x"FA", x"F9", x"FF", x"60", x"F0", x"F0", x"66", x"EF", x"4F", x"06", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"03", x"03", x"00", x"7E", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7E", x"7F", x"7F", x"7F", x"7F", x"BF", x"BF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"80", x"80", x"80", x"80", x"C0", x"C0", x"01", x"01", x"03", x"03", x"03", x"03", x"07", x"07", x"03", x"03", x"07", x"07", x"07", x"07", x"0F", x"0F", 
															x"FD", x"FD", x"FD", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BF", x"BF", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"E0", x"E0", x"C0", x"C0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"1F", x"1F", x"0F", x"0F", x"1F", x"1F", x"1F", x"1F", x"3F", x"3F", x"F7", x"F7", x"F7", x"F7", x"F7", x"EF", x"EF", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EF", x"EF", x"EF", x"EF", x"EF", x"F7", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"F8", x"F8", x"F0", x"F0", x"F8", x"F8", x"F8", x"F8", x"FC", x"FC", x"1F", x"1F", x"1F", x"3F", x"3F", x"3F", x"3F", x"7F", x"3F", x"3F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", 
															x"E0", x"CF", x"DF", x"DF", x"DF", x"DF", x"9F", x"BF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"F3", x"FB", x"FB", x"FB", x"FB", x"F9", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"F8", x"F8", x"FC", x"FC", x"FC", x"FC", x"FE", x"FC", x"FC", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"03", x"03", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BF", x"BF", x"BF", x"3F", x"3F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FD", x"FD", x"FD", x"FC", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"C0", x"C0", x"00", x"00", x"7F", x"FF", x"7F", x"7F", x"FF", x"7F", x"FF", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"7F", x"FF", x"7F", x"7F", x"FF", x"7F", x"7F", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"DB", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"E3", x"F3", x"FF", x"FF", x"FF", x"00", x"0C", x"1E", x"1E", x"3C", x"CE", x"F2", x"FC", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"E0", x"04", x"07", x"04", x"04", x"07", x"04", x"07", x"07", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"92", x"FF", x"92", x"92", x"FF", x"92", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4F", x"FF", x"4F", x"4F", x"FF", x"4F", x"FF", x"FF", x"16", x"00", x"16", x"16", x"00", x"36", x"00", x"00", x"FD", x"FF", x"FD", x"FD", x"FF", x"F7", x"FF", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"6D", x"6D", x"00", x"6D", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"B6", x"B6", x"00", x"B6", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", 
															x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"00", x"00", x"BF", x"FF", x"BF", x"FF", x"FF", x"EF", x"FF", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"00", x"00", x"F2", x"FF", x"F2", x"F2", x"FF", x"F2", x"FF", x"FF", x"68", x"00", x"68", x"68", x"00", x"6C", x"00", x"00", x"49", x"FF", x"49", x"49", x"FF", x"49", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"07", x"20", x"E0", x"20", x"20", x"E0", x"20", x"E0", x"E0", x"07", x"07", x"07", x"07", x"07", x"07", x"04", x"07", x"04", x"04", x"07", x"04", x"04", x"07", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"92", x"FF", x"92", x"92", x"FF", x"92", x"92", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5F", x"FF", x"5F", x"5F", x"FF", x"7F", x"7F", x"FF", x"36", x"00", x"36", x"36", x"00", x"36", x"B6", x"00", 
															x"F7", x"FF", x"F7", x"F7", x"FF", x"E7", x"E7", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"DB", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"6D", x"6D", x"00", x"6D", x"6D", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"B6", x"B6", x"00", x"B6", x"B6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"DB", x"00", x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"DB", x"00", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C3", x"83", x"FF", x"FE", x"FC", x"F8", x"F0", x"E7", x"C4", x"84", x"EF", x"FF", x"EF", x"EF", x"FF", x"E7", x"E7", x"FF", x"DB", x"00", x"DB", x"DB", x"00", x"DB", x"DB", x"00", x"F2", x"FF", x"FA", x"FA", x"FF", x"FE", x"FE", x"FF", x"6C", x"00", x"6C", x"6C", x"00", x"6C", x"6D", x"00", 
															x"49", x"FF", x"49", x"49", x"FF", x"49", x"49", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"E0", x"20", x"20", x"E0", x"20", x"20", x"E0", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"C0", x"40", x"40", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", 
															x"CC", x"C4", x"C4", x"C0", x"C8", x"C8", x"CC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"9F", x"F4", x"92", x"92", x"92", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"C3", x"66", x"66", x"66", x"67", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1A", x"49", x"09", x"79", x"19", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"70", x"24", x"24", x"24", x"30", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C7", x"93", x"93", x"93", x"C7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"03", x"0F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"C0", x"F0", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", x"00", x"00", x"01", x"07", x"0F", x"07", x"01", x"00", x"00", x"03", x"01", x"07", x"0E", x"00", x"01", x"00", x"00", x"00", x"01", x"03", x"07", x"03", x"01", x"00", x"00", x"03", x"01", x"03", x"06", x"00", x"01", x"00", x"00", x"00", x"F8", x"F8", x"F8", x"FC", x"F0", x"78", x"F0", x"F8", x"00", x"40", x"C0", x"C0", x"F0", x"80", 
															x"00", x"00", x"01", x"01", x"03", x"03", x"01", x"00", x"00", x"03", x"01", x"00", x"03", x"00", x"01", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"78", x"F8", x"FC", x"F0", x"B4", x"DC", x"0C", x"F8", x"80", x"FF", x"A0", x"40", x"60", x"60", x"B0", x"C0", x"F8", x"00", x"5F", x"BF", x"9F", x"9F", x"4F", x"3F", x"07", x"FF", x"0B", x"25", x"2D", x"4D", x"5B", x"87", x"3F", x"00", x"F4", x"FA", x"F2", x"F2", x"E4", x"F8", x"C0", x"FE", x"FE", x"FC", x"F0", x"F0", x"F0", x"F0", x"F0", x"01", x"01", x"03", x"0F", x"00", x"00", x"00", x"00", x"FF", x"FF", x"7F", x"1F", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"80", x"E0", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"EF", x"CF", x"CF", x"CF", x"DF", x"DF", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F3", x"F3", x"F3", x"FB", x"FB", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"01", x"01", x"01", x"01", x"03", x"03", x"9F", x"BF", x"BF", x"3F", x"3F", x"3F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F9", x"FD", x"FD", x"FC", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"1F", x"1F", x"1F", x"1F", x"3F", x"3F", x"3F", x"3F", x"3F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", 
															x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"F8", x"F8", x"F8", x"F8", x"FC", x"FC", x"FC", x"FC", x"FC", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"03", x"03", x"3F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FD", x"FD", x"F9", x"F9", x"F9", x"FB", x"FB", x"F3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"BF", x"BF", x"9F", x"9F", x"9F", x"DF", x"DF", x"CF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"C0", x"C0", x"00", x"01", x"01", x"01", x"01", x"03", x"03", x"03", x"03", x"03", x"07", x"07", x"07", x"07", x"0F", x"0F", x"F3", x"F3", x"F7", x"F7", x"E7", x"E7", x"E7", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CF", x"CF", x"EF", x"EF", x"E7", x"E7", x"E7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"80", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"03", x"07", x"07", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"1F", x"3F", x"3F", 
															x"EF", x"CF", x"CF", x"CF", x"DF", x"DF", x"9F", x"9F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F3", x"F3", x"F3", x"FB", x"FB", x"F9", x"F9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F8", x"F8", x"F8", x"F8", x"FC", x"FC", x"0F", x"1F", x"1F", x"1F", x"1F", x"3F", x"00", x"00", x"3F", x"3F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"BF", x"BF", x"3F", x"3F", x"3F", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"F9", x"FD", x"FD", x"FC", x"FC", x"FC", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"F8", x"F8", x"F8", x"F8", x"FC", x"00", x"00", x"FC", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"07", x"17", x"1E", x"0C", x"00", x"00", x"01", x"01", x"00", x"00", x"05", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"05", x"0D", x"0B", x"0A", x"0F", x"1A", x"17", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"14", x"14", x"34", x"2C", x"28", x"3F", x"68", x"5F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"50", x"50", x"D0", x"B0", x"90", x"B0", x"20", x"20", x"00", x"3F", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"FF", x"C0", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"00", x"00", x"F8", x"FC", x"FC", x"FC", x"F0", x"78", x"F0", x"F8", x"C0", x"68", x"C8", x"70", x"F0", x"80", 
															x"98", x"78", x"F8", x"80", x"38", x"70", x"00", x"00", x"62", x"82", x"C2", x"FE", x"C4", x"84", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"14", x"14", x"14", x"14", x"14", x"F4", x"1C", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0A", x"0A", x"0A", x"0A", x"0A", x"FA", x"0E", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"09", x"09", x"09", x"09", x"09", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"1F", x"1F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FF", x"FF", x"3F", x"1F", x"0F", x"07", x"07", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"FF", x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"81", x"00", x"63", x"73", x"7B", x"7F", x"6F", x"67", x"63", x"FF", x"9C", x"8C", x"84", x"80", x"90", x"98", x"9C", x"00", x"0C", x"0C", x"0C", x"08", x"00", x"18", x"18", x"FF", x"F3", x"F3", x"F3", x"F7", x"FF", x"E7", x"E7", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"1F", x"1F", x"0F", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1F", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"F8", x"F8", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"38", x"18", x"0C", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"66", x"66", x"66", x"3C", x"FF", x"C3", x"99", x"99", x"99", x"99", x"99", x"C3", x"00", x"66", x"66", x"66", x"66", x"66", x"66", x"3C", x"FF", x"99", x"99", x"99", x"99", x"99", x"99", x"C3", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"FF", x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"00", x"3F", x"30", x"30", x"3F", x"30", x"30", x"3F", x"FF", x"C0", x"CF", x"CF", x"C0", x"CF", x"CF", x"C0", x"00", x"F8", x"C1", x"C3", x"F3", x"C3", x"C3", x"C3", x"FF", x"07", x"3E", x"3C", x"0C", x"3C", x"3C", x"3C", 
															x"00", x"C6", x"E6", x"36", x"36", x"F6", x"36", x"33", x"FF", x"39", x"19", x"C9", x"C9", x"09", x"C9", x"CC", x"00", x"66", x"66", x"66", x"66", x"66", x"66", x"C7", x"FF", x"99", x"99", x"99", x"99", x"99", x"99", x"38", x"00", x"3F", x"0C", x"0C", x"0C", x"0C", x"0C", x"CC", x"FF", x"C0", x"F3", x"F3", x"F3", x"F3", x"F3", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"78", x"38", x"38", x"18", x"0C", x"00", x"00", x"F8", x"CD", x"CD", x"CD", x"CD", x"CD", x"F8", x"00", x"07", x"32", x"32", x"32", x"32", x"32", x"07", x"FF", x"F3", x"9B", x"9B", x"9B", x"9B", x"9B", x"F1", x"00", x"0C", x"64", x"64", x"64", x"64", x"64", x"0E", x"FF", x"37", x"36", x"36", x"37", x"36", x"36", x"E7", x"00", x"C8", x"C9", x"C9", x"C8", x"C9", x"C9", x"18", x"FF", x"CC", x"6C", x"6C", x"CC", x"6C", x"6C", x"CF", x"00", x"33", x"93", x"93", x"33", x"93", x"93", x"30", x"FF", 
															x"3E", x"30", x"30", x"3E", x"30", x"30", x"BE", x"00", x"C1", x"CF", x"CF", x"C1", x"CF", x"CF", x"41", x"FF", x"00", x"FB", x"C3", x"C3", x"FB", x"C3", x"C3", x"F9", x"FF", x"04", x"3C", x"3C", x"04", x"3C", x"3C", x"06", x"00", x"33", x"36", x"36", x"36", x"36", x"36", x"E3", x"FF", x"CC", x"C9", x"C9", x"C9", x"C9", x"C9", x"1C", x"00", x"CF", x"6C", x"0C", x"0F", x"0C", x"6C", x"CF", x"FF", x"30", x"93", x"F3", x"F0", x"F3", x"93", x"30", x"00", x"86", x"06", x"06", x"84", x"00", x"0C", x"8C", x"FF", x"79", x"F9", x"F9", x"7B", x"FF", x"F3", x"73", x"00", x"7C", x"66", x"66", x"66", x"66", x"66", x"7C", x"FF", x"83", x"99", x"99", x"99", x"99", x"99", x"83", x"03", x"07", x"07", x"0F", x"0F", x"07", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"EF", x"C7", x"03", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FD", 
															x"FF", x"80", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"80", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C0", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E0", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
															x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"08", x"0F", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"00", x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"10", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BC", x"BD", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"BD", x"BD", x"BD", x"BD", x"BD", x"BD", x"BD", x"BD", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"BD", x"BC", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"7E", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"80", x"BE", x"BE", x"BF", x"BF", x"BF", x"BF", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", 
															x"00", x"80", x"80", x"40", x"20", x"A0", x"90", x"C8", x"00", x"00", x"00", x"80", x"C0", x"C0", x"E0", x"F0", x"FF", x"81", x"BD", x"BD", x"BD", x"BD", x"BD", x"BD", x"00", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"E8", x"E4", x"F2", x"FA", x"F9", x"FC", x"FE", x"FE", x"F0", x"F8", x"FC", x"FC", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"20", x"A0", x"90", x"C8", x"E8", x"E4", x"F2", x"FA", x"C0", x"C0", x"E0", x"F0", x"F0", x"F8", x"FC", x"FC", x"BF", x"BF", x"BF", x"BD", x"BC", x"BC", x"BC", x"BD", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"F9", x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BD", x"BD", x"BD", x"3D", x"3D", x"BD", x"BD", x"FD", x"7E", x"7E", x"7E", x"FE", x"FE", x"FE", x"FE", x"FE", x"BF", x"9F", x"4F", x"2F", x"27", x"13", x"0B", x"09", x"7F", x"7F", x"3F", x"1F", x"1F", x"0F", x"07", x"07", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"04", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"7F", x"3F", x"BF", x"9F", x"4F", x"2F", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"3F", x"1F", x"27", x"13", x"0B", x"09", x"04", x"02", x"02", x"01", x"1F", x"0F", x"07", x"07", x"03", x"01", x"01", x"00", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"7D", x"3D", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", 
															x"01", x"02", x"04", x"09", x"13", x"27", x"4F", x"9F", x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"80", x"40", x"20", x"90", x"C8", x"E4", x"F2", x"F9", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"9F", x"4F", x"27", x"13", x"09", x"04", x"02", x"01", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", x"00", x"F9", x"F2", x"E4", x"C8", x"90", x"20", x"40", x"80", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"00", x"BD", x"BD", x"BD", x"BD", x"BD", x"BD", x"81", x"FF", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"00", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"3D", x"BD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"7E", x"BD", x"3D", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"7E", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"97", x"83", x"AB", x"AB", x"AB", x"FF", x"00", x"00", x"68", x"7C", x"54", x"54", x"54", x"00");
	
	constant EXCITEBIKE_CHR_ROM : CHR_ROM_ARRAY := (x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"01", x"0C", x"18", x"30", x"24", x"27", x"31", x"1B", x"0E", x"0F", x"1B", x"33", x"24", x"20", x"31", x"1B", x"0E", x"00", x"00", x"00", x"3C", x"7C", x"78", x"0E", x"7E", x"00", x"00", x"00", x"00", x"02", x"07", x"7E", x"04", x"4F", x"C0", x"C8", x"C0", x"E2", x"E3", x"F1", x"F9", x"70", x"38", x"70", x"BE", x"9F", x"C0", x"66", x"A6", x"78", x"78", x"45", x"C5", x"81", x"81", x"08", x"00", x"D7", x"C6", x"3D", x"3D", x"39", x"BD", x"08", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"00", x"80", x"00", x"00", x"00", x"80", x"80", x"80", x"F0", x"08", 
															x"F0", x"D8", x"CC", x"64", x"24", x"8C", x"D8", x"70", x"30", x"18", x"8C", x"04", x"04", x"8C", x"D8", x"70", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"08", x"10", x"14", x"10", x"19", x"0F", x"0F", x"07", x"0B", x"13", x"13", x"10", x"19", x"0F", x"00", x"00", x"00", x"3C", x"7C", x"78", x"0E", x"7E", x"00", x"00", x"00", x"00", x"02", x"07", x"7E", x"04", x"4F", x"C0", x"C8", x"C8", x"C0", x"E0", x"F2", x"7B", x"70", x"38", x"70", x"B0", x"B8", x"DE", x"6F", x"20", x"F9", x"F9", x"44", x"44", x"C5", x"41", x"89", x"00", x"D6", x"C6", x"FF", x"BE", x"3D", x"7D", x"89", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"00", x"E0", x"D0", x"E8", x"64", x"04", x"8C", x"F0", x"F0", x"28", x"10", x"88", x"04", x"04", x"8C", x"F0", 
															x"00", x"00", x"00", x"01", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"0F", x"13", x"0C", x"18", x"31", x"27", x"26", x"31", x"1B", x"0E", x"0F", x"1B", x"31", x"24", x"20", x"31", x"1B", x"0E", x"00", x"00", x"F0", x"F0", x"E0", x"38", x"F8", x"3C", x"00", x"00", x"00", x"08", x"1C", x"F8", x"10", x"C0", x"00", x"01", x"85", x"C7", x"E3", x"F1", x"F1", x"79", x"E0", x"FD", x"7F", x"01", x"8C", x"4E", x"2E", x"D7", x"71", x"C1", x"81", x"80", x"88", x"80", x"00", x"00", x"C9", x"79", x"39", x"3C", x"98", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"D8", x"8C", x"00", x"00", x"00", x"E0", x"00", x"70", x"58", x"0C", x"E4", x"A4", x"8C", x"D8", x"70", x"00", x"00", x"00", x"04", x"84", x"8C", x"D8", x"70", x"00", x"00", x"00", 
															x"00", x"07", x"0F", x"0F", x"01", x"0F", x"09", x"08", x"00", x"00", x"00", x"00", x"0F", x"00", x"0E", x"07", x"08", x"0C", x"0F", x"0F", x"07", x"07", x"07", x"0D", x"07", x"07", x"06", x"02", x"03", x"00", x"07", x"3F", x"00", x"11", x"31", x"21", x"27", x"31", x"1B", x"0E", x"0E", x"1F", x"36", x"20", x"24", x"31", x"1B", x"0E", x"00", x"80", x"80", x"00", x"C0", x"C0", x"E8", x"88", x"00", x"00", x"40", x"E0", x"C0", x"80", x"08", x"89", x"14", x"08", x"0F", x"C3", x"E3", x"F3", x"E3", x"81", x"FF", x"E4", x"11", x"1C", x"9E", x"5A", x"13", x"71", x"00", x"80", x"88", x"80", x"80", x"80", x"00", x"00", x"F8", x"7C", x"38", x"80", x"80", x"80", x"00", x"00", x"00", x"E0", x"B0", x"18", x"08", x"C8", x"18", x"B0", x"00", x"E0", x"B0", x"18", x"08", x"08", x"18", x"B0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"03", x"07", x"07", x"00", x"07", x"04", x"0C", x"0C", x"00", x"00", x"00", x"07", x"00", x"07", x"03", x"03", x"0C", x"0E", x"0F", x"0F", x"07", x"03", x"06", x"00", x"07", x"05", x"04", x"03", x"00", x"03", x"0F", x"0B", x"00", x"04", x"0C", x"08", x"09", x"0C", x"06", x"03", x"13", x"07", x"0C", x"08", x"09", x"0C", x"06", x"03", x"C0", x"C0", x"80", x"E0", x"E0", x"F8", x"88", x"14", x"00", x"20", x"70", x"E0", x"40", x"08", x"89", x"FF", x"0D", x"07", x"E2", x"F2", x"FB", x"E1", x"40", x"40", x"E3", x"98", x"3E", x"8E", x"6B", x"19", x"FC", x"FE", x"60", x"E4", x"60", x"E0", x"A0", x"60", x"C0", x"80", x"DF", x"8C", x"20", x"20", x"20", x"60", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"E0", x"B0", x"98", x"C8", x"48", x"18", x"B0", x"E0", x"00", x"B0", x"18", x"08", x"08", x"18", x"B0", x"E0", x"00", 
															x"0F", x"1F", x"1E", x"03", x"1F", x"13", x"32", x"30", x"00", x"00", x"01", x"1F", x"01", x"1C", x"0E", x"0F", x"30", x"39", x"1F", x"0F", x"01", x"03", x"03", x"02", x"1F", x"0E", x"07", x"00", x"00", x"03", x"03", x"07", x"00", x"00", x"03", x"02", x"02", x"03", x"01", x"00", x"0D", x"09", x"13", x"02", x"02", x"03", x"01", x"00", x"00", x"00", x"00", x"80", x"A1", x"F3", x"1F", x"4F", x"00", x"80", x"C2", x"84", x"25", x"3B", x"20", x"C0", x"03", x"C1", x"F0", x"EC", x"E4", x"C0", x"C4", x"30", x"9B", x"3D", x"18", x"DC", x"1E", x"BE", x"FC", x"E8", x"30", x"30", x"38", x"28", x"68", x"18", x"B0", x"E0", x"C0", x"90", x"98", x"08", x"48", x"18", x"B0", x"E0", x"00", x"00", x"00", x"E0", x"B0", x"18", x"08", x"C8", x"00", x"00", x"00", x"E0", x"B0", x"18", x"08", x"08", x"18", x"B0", x"E0", x"00", x"00", x"00", x"00", x"00", x"18", x"B0", x"E0", x"00", x"00", x"00", x"00", x"00", 
															x"1E", x"3E", x"3C", x"07", x"3F", x"27", x"62", x"60", x"00", x"01", x"03", x"3F", x"02", x"38", x"1E", x"3C", x"70", x"30", x"3F", x"1F", x"1F", x"0F", x"03", x"03", x"1F", x"0F", x"09", x"0E", x"00", x"01", x"03", x"03", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"05", x"05", x"0D", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"21", x"93", x"1F", x"32", x"00", x"00", x"82", x"06", x"25", x"1B", x"20", x"E2", x"03", x"61", x"F8", x"F4", x"E0", x"C0", x"A0", x"34", x"DF", x"9D", x"4C", x"0C", x"DC", x"FE", x"FF", x"CC", x"30", x"18", x"1C", x"14", x"14", x"8C", x"D8", x"70", x"E0", x"C8", x"8C", x"04", x"04", x"8C", x"D8", x"70", x"00", x"00", x"00", x"E0", x"B0", x"18", x"C8", x"48", x"00", x"00", x"00", x"E0", x"B0", x"18", x"08", x"08", x"18", x"B0", x"E0", x"00", x"00", x"00", x"00", x"00", x"18", x"B0", x"E0", x"00", x"00", x"00", x"00", x"00", 
															x"07", x"0F", x"0F", x"01", x"0F", x"09", x"18", x"18", x"00", x"00", x"00", x"0F", x"00", x"0E", x"07", x"07", x"18", x"1C", x"1E", x"0F", x"0F", x"07", x"03", x"00", x"07", x"07", x"05", x"06", x"01", x"00", x"00", x"00", x"80", x"80", x"01", x"C3", x"C2", x"E3", x"83", x"3F", x"00", x"40", x"E1", x"CB", x"8A", x"08", x"89", x"B1", x"08", x"10", x"1B", x"FC", x"F8", x"F8", x"CE", x"0D", x"14", x"FF", x"E7", x"33", x"C7", x"07", x"0F", x"0E", x"0C", x"0C", x"00", x"02", x"02", x"03", x"01", x"00", x"0F", x"0F", x"0B", x"0A", x"0A", x"0B", x"01", x"00", x"00", x"E0", x"B0", x"18", x"C8", x"C8", x"18", x"B0", x"00", x"E0", x"B0", x"18", x"08", x"08", x"18", x"B0", x"E0", x"00", x"C0", x"00", x"00", x"40", x"00", x"80", x"E0", x"00", x"C0", x"E0", x"C0", x"C0", x"80", x"00", x"E0", x"F0", x"58", x"48", x"48", x"18", x"B0", x"E0", x"20", x"30", x"18", x"08", x"08", x"18", x"B0", x"E0", 
															x"07", x"0D", x"18", x"13", x"11", x"19", x"0D", x"07", x"07", x"0D", x"18", x"10", x"10", x"18", x"0C", x"06", x"01", x"01", x"03", x"03", x"04", x"00", x"00", x"00", x"08", x"06", x"02", x"02", x"05", x"00", x"00", x"00", x"00", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"01", x"00", x"00", x"00", x"80", x"C0", x"40", x"40", x"C4", x"80", x"20", x"00", x"80", x"C0", x"40", x"40", x"DC", x"8C", x"2E", x"21", x"1B", x"3E", x"7C", x"8E", x"07", x"07", x"03", x"FE", x"E4", x"D3", x"53", x"F9", x"FC", x"3C", x"3E", x"03", x"E3", x"FF", x"C6", x"78", x"F8", x"F0", x"00", x"1E", x"3C", x"84", x"F8", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"D8", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"D8", x"8C", x"E4", x"04", x"0C", x"18", x"70", x"80", x"80", x"0C", x"04", x"84", x"CC", x"D8", x"F0", x"00", x"70", 
															x"0E", x"1B", x"31", x"24", x"24", x"37", x"1B", x"0F", x"0E", x"1B", x"31", x"20", x"20", x"31", x"19", x"0C", x"01", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"0F", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"07", x"03", x"03", x"00", x"01", x"01", x"00", x"00", x"00", x"01", x"03", x"07", x"02", x"00", x"00", x"00", x"10", x"81", x"81", x"A3", x"A3", x"1E", x"1E", x"00", x"10", x"BD", x"9C", x"BC", x"BD", x"63", x"EB", x"9D", x"8F", x"CF", x"4F", x"07", x"07", x"03", x"03", x"65", x"66", x"03", x"F1", x"79", x"3A", x"1E", x"1E", x"43", x"C3", x"FE", x"80", x"F0", x"F0", x"E0", x"00", x"7E", x"7C", x"08", x"F0", x"00", x"00", x"00", x"00", x"70", x"D8", x"8C", x"E4", x"24", x"0C", x"18", x"30", x"70", x"D8", x"8C", x"04", x"24", x"CC", x"D8", x"F0", x"80", x"80", x"80", x"F0", x"F0", x"F0", x"E0", x"C0", x"80", x"70", x"00", x"09", x"7F", x"4F", x"8E", x"00", 
															x"00", x"07", x"0D", x"18", x"12", x"13", x"19", x"0D", x"00", x"07", x"0D", x"18", x"10", x"10", x"18", x"0D", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"06", x"05", x"07", x"06", x"07", x"06", x"01", x"03", x"06", x"04", x"04", x"04", x"11", x"3B", x"00", x"06", x"8F", x"DF", x"4F", x"47", x"C1", x"F0", x"79", x"7B", x"90", x"D4", x"72", x"79", x"38", x"09", x"14", x"10", x"7E", x"3F", x"38", x"0F", x"1F", x"1E", x"67", x"9F", x"0F", x"10", x"3F", x"70", x"20", x"00", x"C0", x"60", x"30", x"90", x"10", x"30", x"20", x"00", x"C0", x"60", x"30", x"90", x"10", x"30", x"E0", x"D9", x"40", x"C0", x"C0", x"80", x"DC", x"FE", x"FE", x"78", x"F3", x"E7", x"C7", x"8F", x"02", x"88", x"50", x"C0", x"38", x"0C", x"0C", x"1C", x"BC", x"F0", x"C0", x"00", x"F0", x"F0", x"F0", x"F8", x"C0", x"80", x"80", x"00", 
															x"07", x"0D", x"18", x"12", x"16", x"1A", x"0F", x"07", x"07", x"0D", x"18", x"10", x"10", x"18", x"0C", x"04", x"01", x"00", x"00", x"04", x"00", x"00", x"00", x"07", x"00", x"01", x"03", x"07", x"03", x"02", x"00", x"07", x"0D", x"18", x"13", x"13", x"18", x"0D", x"07", x"00", x"0D", x"18", x"10", x"10", x"18", x"0D", x"07", x"00", x"00", x"80", x"C0", x"40", x"00", x"80", x"99", x"19", x"00", x"80", x"C1", x"48", x"68", x"E8", x"F8", x"78", x"59", x"39", x"1F", x"1F", x"3F", x"DC", x"04", x"18", x"78", x"C0", x"E0", x"E8", x"C7", x"E3", x"F7", x"44", x"FE", x"E0", x"C3", x"41", x"C0", x"80", x"00", x"00", x"8E", x"88", x"08", x"48", x"C8", x"83", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"00", x"00", x"E0", x"E0", x"E0", x"E0", x"00", x"80", x"C0", x"C0", x"E0", x"F8", x"FC", x"0E", x"0E", x"06", x"80", x"80", x"40", x"00", x"90", x"F8", x"F8", x"78", 
															x"06", x"06", x"CC", x"F8", x"C0", x"78", x"F8", x"F0", x"F8", x"78", x"38", x"80", x"F8", x"80", x"00", x"00", x"00", x"00", x"01", x"03", x"06", x"04", x"04", x"06", x"00", x"00", x"01", x"03", x"06", x"04", x"04", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C3", x"63", x"37", x"8F", x"86", x"E6", x"00", x"00", x"C8", x"68", x"38", x"93", x"39", x"3D", x"66", x"FE", x"17", x"07", x"02", x"02", x"20", x"00", x"3D", x"89", x"1A", x"18", x"3C", x"3F", x"31", x"10", x"03", x"06", x"0C", x"09", x"09", x"0C", x"06", x"03", x"03", x"06", x"0C", x"08", x"08", x"0C", x"06", x"03", x"3C", x"7C", x"F8", x"8E", x"FE", x"1F", x"00", x"00", x"00", x"02", x"87", x"FE", x"84", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"A0", x"00", x"18", x"50", x"40", x"80", x"E0", x"E0", x"E0", x"90", x"D8", x"B0", x"20", 
															x"C0", x"C0", x"E0", x"A0", x"20", x"60", x"C0", x"80", x"10", x"50", x"60", x"20", x"20", x"60", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"1C", x"36", x"63", x"00", x"00", x"00", x"00", x"01", x"1C", x"36", x"63", x"40", x"48", x"6F", x"37", x"1C", x"00", x"00", x"00", x"41", x"49", x"61", x"34", x"1C", x"00", x"00", x"00", x"00", x"01", x"03", x"1F", x"3C", x"73", x"60", x"60", x"00", x"00", x"00", x"04", x"07", x"9C", x"1F", x"9C", x"70", x"38", x"3D", x"FC", x"C9", x"45", x"05", x"49", x"DE", x"CF", x"CB", x"50", x"36", x"7E", x"7E", x"78", x"03", x"07", x"0D", x"09", x"09", x"0C", x"06", x"03", x"32", x"16", x"0C", x"08", x"08", x"0C", x"06", x"03", x"00", x"E0", x"E0", x"C0", x"70", x"F0", x"F8", x"00", x"00", x"00", x"10", x"38", x"F0", x"20", x"80", x"00", x"00", x"00", x"40", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"40", x"80", x"80", x"80", x"C0", x"60", 
															x"80", x"C0", x"60", x"20", x"20", x"60", x"C0", x"80", x"80", x"C0", x"60", x"20", x"20", x"60", x"C0", x"80", x"0E", x"1A", x"30", x"24", x"27", x"31", x"1B", x"0E", x"0F", x"1B", x"31", x"24", x"20", x"30", x"1B", x"0E", x"00", x"03", x"07", x"3F", x"78", x"77", x"60", x"60", x"00", x"00", x"00", x"08", x"0F", x"B8", x"BF", x"9E", x"E0", x"30", x"38", x"7C", x"DD", x"88", x"80", x"40", x"DC", x"CF", x"EF", x"C9", x"E3", x"77", x"7A", x"7B", x"01", x"03", x"07", x"05", x"05", x"06", x"03", x"01", x"33", x"12", x"06", x"04", x"04", x"06", x"03", x"01", x"00", x"C0", x"C0", x"80", x"E0", x"E0", x"F0", x"00", x"00", x"00", x"20", x"70", x"E0", x"40", x"00", x"00", x"00", x"00", x"00", x"B0", x"A0", x"80", x"80", x"80", x"00", x"00", x"80", x"B0", x"60", x"00", x"40", x"30", x"C0", x"E0", x"30", x"90", x"90", x"30", x"60", x"C0", x"50", x"60", x"30", x"10", x"10", x"30", x"60", x"C0", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"0E", x"18", x"30", x"24", x"27", x"0C", x"06", x"01", x"0F", x"1B", x"33", x"25", x"20", x"31", x"1B", x"0E", x"00", x"00", x"00", x"00", x"00", x"31", x"1B", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"1E", x"63", x"FF", x"C7", x"C0", x"00", x"00", x"00", x"01", x"3F", x"21", x"7C", x"38", x"C0", x"E0", x"E0", x"F1", x"7C", x"5C", x"4C", x"84", x"BC", x"7C", x"1F", x"CF", x"D8", x"E3", x"F7", x"7F", x"8D", x"01", x"23", x"02", x"02", x"03", x"01", x"00", x"7F", x"31", x"3B", x"02", x"02", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"00", x"00", x"00", x"80", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"C0", x"C0", x"80", x"80", x"00", x"00", x"00", x"A0", x"40", x"40", x"60", x"10", 
															x"E0", x"B0", x"98", x"88", x"C8", x"18", x"B0", x"E0", x"60", x"30", x"18", x"08", x"08", x"18", x"B0", x"E0", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"00", x"00", x"07", x"03", x"03", x"00", x"78", x"38", x"3A", x"01", x"3C", x"61", x"4F", x"7F", x"7F", x"3F", x"00", x"3E", x"7F", x"62", x"40", x"7F", x"7F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"04", x"03", x"07", x"C1", x"C3", x"E3", x"00", x"00", x"83", x"C4", x"C0", x"1E", x"9F", x"9C", x"FE", x"71", x"FC", x"FC", x"FD", x"BD", x"9D", x"00", x"C3", x"FE", x"07", x"3E", x"BD", x"BD", x"9D", x"00", x"00", x"C0", x"80", x"40", x"E0", x"1C", x"36", x"E6", x"00", x"00", x"60", x"F8", x"F8", x"FC", x"F6", x"A6", x"6E", x"FC", x"FC", x"9C", x"B8", x"F8", x"F0", x"E0", x"EE", x"1C", x"DC", x"9C", x"B8", x"F8", x"F0", x"E0", 
															x"00", x"01", x"02", x"02", x"03", x"03", x"03", x"01", x"00", x"00", x"01", x"01", x"00", x"10", x"3F", x"3F", x"1E", x"30", x"61", x"4F", x"63", x"7F", x"3E", x"00", x"3F", x"33", x"60", x"40", x"63", x"7F", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BF", x"38", x"3F", x"0F", x"06", x"80", x"F2", x"FB", x"50", x"CF", x"E7", x"C0", x"F4", x"7D", x"1C", x"C0", x"61", x"63", x"FE", x"FE", x"3C", x"1C", x"04", x"00", x"FE", x"FF", x"1A", x"77", x"EF", x"FC", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B8", x"6C", x"80", x"80", x"00", x"18", x"3C", x"78", x"78", x"EC", x"CC", x"EC", x"AC", x"9C", x"98", x"B8", x"F0", x"60", x"4C", x"0C", x"8C", x"9C", x"98", x"B8", x"F0", x"60", x"00", x"00", x"19", x"7F", x"7F", x"1F", x"0F", x"01", x"F0", x"70", x"60", x"10", x"0B", x"04", x"00", x"1F", 
															x"00", x"1C", x"30", x"65", x"4F", x"61", x"3F", x"1E", x"03", x"1F", x"33", x"67", x"40", x"61", x"3F", x"1E", x"00", x"00", x"00", x"07", x"0F", x"0F", x"01", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"00", x"44", x"C0", x"C0", x"F2", x"F9", x"C1", x"E0", x"F0", x"3C", x"3C", x"7E", x"8E", x"01", x"00", x"03", x"87", x"60", x"74", x"FD", x"FD", x"BD", x"BD", x"01", x"00", x"FF", x"8F", x"05", x"3D", x"FD", x"FD", x"E1", x"70", x"00", x"00", x"00", x"80", x"80", x"00", x"C0", x"80", x"00", x"00", x"00", x"00", x"40", x"E0", x"C0", x"80", x"E0", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"78", x"C0", x"F8", x"EC", x"24", x"24", x"8C", x"FC", x"F8", x"08", x"B8", x"8C", x"04", x"04", x"8C", x"FC", x"F8", x"00", x"01", x"01", x"01", x"03", x"03", x"23", x"73", x"00", x"00", x"00", x"00", x"02", x"1E", x"3E", x"7F", 
															x"7C", x"60", x"6F", x"23", x"1E", x"00", x"00", x"00", x"7F", x"63", x"60", x"20", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"41", x"2E", x"E0", x"3F", x"1E", x"1C", x"08", x"87", x"C1", x"FB", x"7F", x"DF", x"E1", x"F0", x"E8", x"FF", x"BC", x"4E", x"F6", x"76", x"8C", x"8C", x"00", x"00", x"00", x"00", x"4E", x"0E", x"7F", x"7C", x"70", x"38", x"00", x"00", x"80", x"00", x"00", x"20", x"40", x"C0", x"E0", x"A0", x"00", x"C0", x"F0", x"70", x"40", x"C0", x"C0", x"80", x"80", x"E0", x"58", x"6C", x"6C", x"4C", x"2C", x"18", x"78", x"3C", x"18", x"0C", x"4C", x"4C", x"2C", x"18", x"00", x"01", x"01", x"01", x"01", x"03", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"02", x"0F", x"1F", x"00", x"0E", x"18", x"19", x"1B", x"18", x"1F", x"0F", x"1F", x"0F", x"19", x"18", x"18", x"18", x"1F", x"0F", 
															x"00", x"00", x"00", x"3E", x"7E", x"63", x"5F", x"26", x"00", x"00", x"00", x"00", x"01", x"1F", x"21", x"59", x"C0", x"C0", x"F1", x"FB", x"F9", x"FD", x"FC", x"9C", x"3F", x"3F", x"0F", x"42", x"46", x"72", x"0B", x"E3", x"32", x"22", x"62", x"A0", x"88", x"88", x"80", x"00", x"EF", x"DE", x"BE", x"3E", x"9E", x"88", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"E0", x"20", x"C0", x"80", x"80", x"80", x"80", x"B0", x"D0", x"E0", x"C0", x"80", x"80", x"00", x"70", x"78", x"10", x"E8", x"A8", x"88", x"98", x"D0", x"60", x"00", x"00", x"88", x"88", x"88", x"98", x"D0", x"60", x"00", x"00", x"78", x"78", x"C5", x"C5", x"C1", x"81", x"28", x"00", x"D7", x"C6", x"BD", x"3D", x"79", x"FD", x"E8", x"70", x"00", x"00", x"78", x"E1", x"C1", x"3F", x"F7", x"62", x"01", x"01", x"01", x"1C", x"3E", x"3C", x"1C", x"7C", 
															x"9C", x"88", x"80", x"C1", x"63", x"7F", x"3F", x"1E", x"73", x"77", x"7F", x"3E", x"3E", x"18", x"01", x"03", x"00", x"00", x"00", x"80", x"A1", x"BB", x"1F", x"4F", x"00", x"C0", x"C2", x"04", x"25", x"3F", x"20", x"C0", x"00", x"C0", x"F8", x"EC", x"E4", x"40", x"04", x"30", x"9C", x"3C", x"98", x"5C", x"1E", x"3E", x"3C", x"68", x"00", x"01", x"3C", x"61", x"4F", x"7F", x"7F", x"3F", x"00", x"3E", x"7F", x"62", x"40", x"7F", x"7F", x"3F", x"C2", x"71", x"FC", x"FC", x"FD", x"BD", x"9D", x"00", x"C3", x"FE", x"07", x"3E", x"BD", x"BD", x"9D", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"36", x"A6", x"00", x"00", x"00", x"00", x"00", x"7C", x"F6", x"E6", x"6E", x"FC", x"FC", x"9C", x"B8", x"F8", x"F0", x"E0", x"EE", x"1C", x"DC", x"9C", x"B8", x"F8", x"F0", x"E0", x"81", x"C3", x"81", x"B9", x"BD", x"FB", x"D7", x"82", x"00", x"38", x"BD", x"A9", x"A1", x"C3", x"EF", x"FE", 
															x"38", x"00", x"00", x"7C", x"6C", x"6C", x"00", x"00", x"44", x"7C", x"7C", x"00", x"00", x"00", x"6C", x"EE", x"01", x"03", x"01", x"1D", x"3D", x"1D", x"6B", x"C2", x"00", x"1C", x"3D", x"15", x"05", x"01", x"77", x"FE", x"DC", x"80", x"E0", x"7E", x"36", x"36", x"00", x"00", x"E2", x"BE", x"DE", x"4E", x"36", x"36", x"36", x"77", x"80", x"C1", x"83", x"B9", x"BD", x"FB", x"D7", x"86", x"00", x"38", x"BC", x"A9", x"A1", x"C3", x"EF", x"FE", x"38", x"00", x"00", x"00", x"00", x"6C", x"00", x"00", x"7C", x"7C", x"7C", x"7C", x"6C", x"6C", x"6C", x"EE", x"00", x"00", x"00", x"00", x"FB", x"FD", x"B9", x"D7", x"00", x"00", x"38", x"3C", x"28", x"A0", x"81", x"EF", x"83", x"BA", x"00", x"00", x"00", x"00", x"6C", x"00", x"FF", x"FE", x"7C", x"7C", x"FE", x"C6", x"6C", x"EE", x"3C", x"0E", x"0E", x"70", x"7E", x"7C", x"0E", x"CE", x"00", x"70", x"F0", x"7E", x"51", x"03", x"1D", x"11", 
															x"CF", x"0F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"30", x"78", x"2C", x"00", x"00", x"07", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"80", x"00", x"00", x"00", x"C0", x"E0", x"C0", x"80", x"00", x"C0", x"C0", x"C0", x"C0", x"80", x"00", x"00", x"00", x"80", x"40", x"80", x"80", x"40", x"80", x"C0", x"80", x"3C", x"0E", x"0E", x"70", x"7E", x"7C", x"18", x"18", x"00", x"70", x"F0", x"7E", x"50", x"02", x"3F", x"07", x"68", x"61", x"01", x"3F", x"07", x"03", x"00", x"00", x"17", x"1E", x"3E", x"7A", x"71", x"70", x"F0", x"E0", x"00", x"00", x"80", x"80", x"C0", x"80", x"00", x"00", x"40", x"E0", x"70", x"70", x"10", x"00", x"00", x"00", x"1E", x"8F", x"C6", x"C6", x"40", x"00", x"00", x"00", x"C1", x"FB", x"FF", x"FF", x"63", x"03", x"07", x"07", x"00", x"00", x"1E", x"0F", x"07", x"38", x"3F", x"3E", x"00", x"00", x"00", x"30", x"78", x"3F", x"28", x"01", 
															x"38", x"FC", x"FC", x"7C", x"38", x"36", x"06", x"00", x"FF", x"1F", x"07", x"E7", x"DF", x"C1", x"80", x"80", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EF", x"EF", x"EF", x"C7", x"C7", x"83", x"83", x"01", x"38", x"FE", x"7C", x"00", x"00", x"00", x"00", x"00", x"38", x"FE", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"78", x"3C", x"0E", x"00", x"00", x"00", x"00", x"F0", x"78", x"3C", x"0E", x"00", x"00", x"00", x"00", x"80", x"60", x"70", x"38", x"18", x"0C", x"06", x"00", x"80", x"60", x"70", x"38", x"18", x"0C", x"06", x"60", x"20", x"30", x"10", x"18", x"08", x"0C", x"04", x"60", x"20", x"30", x"10", x"18", x"08", x"0C", x"04", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"06", x"00", x"00", x"06", x"1D", x"1F", x"1F", x"1D", x"01", 
															x"06", x"03", x"03", x"03", x"07", x"0A", x"12", x"20", x"01", x"03", x"00", x"00", x"07", x"0A", x"12", x"20", x"00", x"00", x"1E", x"7E", x"3E", x"24", x"0C", x"3C", x"1E", x"1E", x"03", x"F2", x"F0", x"FE", x"DE", x"DE", x"38", x"1E", x"00", x"00", x"80", x"40", x"20", x"1E", x"DE", x"1E", x"7E", x"7E", x"E6", x"66", x"26", x"1E", x"00", x"00", x"00", x"03", x"43", x"FF", x"FE", x"00", x"00", x"03", x"0F", x"00", x"00", x"3C", x"3F", x"03", x"00", x"00", x"03", x"03", x"07", x"0E", x"0E", x"00", x"03", x"03", x"03", x"03", x"07", x"0E", x"0E", x"1C", x"00", x"00", x"00", x"C0", x"C0", x"E0", x"70", x"30", x"00", x"C0", x"C0", x"00", x"00", x"20", x"F0", x"F0", x"30", x"30", x"F0", x"E0", x"F0", x"70", x"30", x"00", x"F0", x"F0", x"C0", x"E0", x"F0", x"70", x"30", x"38", x"00", x"00", x"1C", x"1C", x"0C", x"1E", x"3E", x"38", x"1C", x"3C", x"00", x"00", x"0C", x"3F", x"77", x"77", 
															x"38", x"3E", x"00", x"00", x"00", x"00", x"00", x"77", x"5F", x"5E", x"3E", x"3E", x"36", x"36", x"36", x"77", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"38", x"38", x"3C", x"26", x"E6", x"EE", x"0C", x"01", x"E1", x"04", x"04", x"3E", x"6E", x"7E", x"72", x"7F", x"E7", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"FF", x"FF", x"7E", x"24", x"24", x"24", x"A5", x"7E", x"FF", x"FF", x"FF", x"DF", x"DF", x"DF", x"5E", 
															x"FF", x"FF", x"FF", x"7E", x"24", x"26", x"24", x"24", x"04", x"04", x"04", x"85", x"DF", x"DD", x"DF", x"5E", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CC", x"CC", x"33", x"33", x"CC", x"CC", x"32", x"32", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"CC", x"CC", x"32", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"01", x"01", x"03", x"03", x"03", x"07", x"00", x"80", x"80", x"80", x"00", x"0F", x"1F", x"0F", x"00", x"00", x"0F", x"4F", x"DF", x"EB", x"63", x"71", x"06", x"08", x"00", x"00", x"3E", x"3E", x"3E", x"00", x"38", x"1E", x"FE", x"FE", x"3E", x"3E", x"3E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8F", x"FE", x"EE", x"EE", x"CE", x"8E", x"8E", x"8E", x"8F", 
															x"00", x"00", x"00", x"00", x"01", x"03", x"01", x"00", x"00", x"01", x"01", x"03", x"01", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"03", x"03", x"03", x"07", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"04", x"03", x"03", x"0C", x"00", x"01", x"01", x"00", x"07", x"03", x"03", x"0C", x"00", x"03", x"03", x"03", x"07", x"00", x"00", x"00", x"00", x"E0", x"E0", x"E0", x"C0", x"00", x"E0", x"E0", x"E0", x"60", x"60", x"20", x"00", x"E0", x"E0", x"70", x"78", x"FC", x"FE", x"FE", x"FF", x"F0", x"F0", x"F0", x"C8", x"30", x"32", x"CC", x"CC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"87", x"33", x"33", x"CC", x"CC", x"33", x"33", x"BC", x"8C", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"08", x"0C", x"0A", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"76", x"49", x"49", x"49", x"45", x"43", x"7F", x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"1C", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2C", x"31", x"31", x"31", x"31", x"2D", x"3F", x"00", x"00", x"20", x"20", x"20", x"20", x"20", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"21", x"21", x"21", x"21", x"21", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"80", x"32", x"0C", x"47", x"09", x"16", x"00", x"08", x"80", x"32", x"0C", x"47", x"09", x"16", x"40", x"AC", x"50", x"18", x"22", x"48", x"32", x"01", x"40", x"AC", x"50", x"18", x"22", x"48", x"32", x"01", 
															x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"40", x"40", x"33", x"33", x"0C", x"0C", x"33", x"33", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1E", x"06", x"06", x"06", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7A", x"43", x"73", x"42", x"7A", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"5C", x"56", x"D2", x"D6", x"5C", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"10", x"10", x"38", x"FE", x"7C", x"38", x"6C", x"44", x"10", x"10", x"38", x"FE", x"7C", x"38", x"6C", x"44", x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F", 
															x"01", x"01", x"01", x"41", x"41", x"41", x"7D", x"39", x"FF", x"E7", x"C3", x"C3", x"C3", x"C3", x"FF", x"FF", x"01", x"01", x"01", x"41", x"41", x"41", x"7D", x"38", x"FF", x"E7", x"C3", x"C3", x"C3", x"C3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"FF", x"FF", x"C3", x"3C", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"3C", x"C3", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C3", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"C3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"00", x"00", x"FF", x"7C", x"38", x"10", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"06", x"38", x"C0", x"00", x"00", x"03", x"02", x"FF", x"F9", x"C7", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"1C", x"03", x"00", x"00", x"C0", x"40", x"FF", x"9F", x"E3", x"FC", x"FF", x"FF", x"FF", x"FF", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"02", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"4E", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"B1", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"36", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"3C", x"99", x"86", x"06", x"00", x"81", x"81", x"C3", x"00", x"60", x"46", x"4E", x"1F", x"9F", x"99", x"89", x"E7", x"C3", x"02", x"18", x"18", x"3C", x"3C", x"3C", x"00", x"00", x"00", x"98", x"D9", x"D9", x"C1", x"81", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"03", x"0C", x"30", x"C0", x"FF", x"FF", x"FF", x"FF", x"FC", x"F3", x"CF", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"F7", x"E7", x"F7", x"F7", x"F7", x"E3", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"E7", x"DB", x"FB", x"E7", x"DF", x"C3", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"33", x"33", x"CC", x"CC", x"33", x"33", x"CC", x"CC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"E7", x"DB", x"F7", x"FB", x"DB", x"E7", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", 
															x"3F", x"3F", x"3F", x"07", x"3B", x"3B", x"39", x"3D", x"C7", x"C7", x"C7", x"FF", x"C7", x"C7", x"C7", x"C7", x"3C", x"3E", x"3E", x"3F", x"3F", x"3F", x"3F", x"3F", x"C7", x"C7", x"C7", x"C7", x"C7", x"C7", x"C7", x"C7", x"7F", x"47", x"47", x"C3", x"83", x"81", x"81", x"81", x"83", x"BB", x"B9", x"3D", x"7C", x"7E", x"7E", x"7E", x"7F", x"80", x"80", x"80", x"80", x"80", x"80", x"7F", x"80", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"80", x"00", x"00", x"00", x"01", x"02", x"04", x"08", x"F0", x"FF", x"FF", x"FF", x"FE", x"FD", x"FB", x"F7", x"0F", x"00", x"00", x"3C", x"3C", x"3C", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", x"00", x"1F", x"1F", x"7F", x"DF", x"9F", x"DF", x"7F", x"00", x"1F", x"11", x"77", x"DF", x"9F", x"DF", x"7F", x"0F", x"07", x"03", x"01", x"03", x"01", x"03", x"07", x"0F", x"07", x"03", x"01", x"03", x"01", x"03", x"07", x"00", x"F8", x"F8", x"FE", x"FB", x"F9", x"FB", x"FE", x"00", x"F8", x"58", x"FE", x"FB", x"F9", x"FB", x"FE", x"F0", x"E0", x"80", x"80", x"C0", x"80", x"C0", x"E0", x"F0", x"E0", x"80", x"80", x"C0", x"80", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", x"00", x"00", x"FF", x"80", x"8F", x"8F", x"8C", x"8C", x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"F3", x"F3", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"8C", x"8E", x"C7", x"63", x"30", x"18", x"0F", x"07", x"F3", x"F1", x"B8", x"9C", x"CF", x"E7", x"F0", x"F8", x"00", x"03", x"07", x"07", x"07", x"07", x"07", x"03", x"FF", x"FC", x"F8", x"F8", x"F8", x"F8", x"F8", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", 
															x"F0", x"F0", x"D0", x"F0", x"F0", x"F0", x"B0", x"F0", x"0F", x"0F", x"2F", x"0F", x"0F", x"0F", x"4F", x"0F", x"F1", x"F1", x"72", x"D2", x"F4", x"F4", x"F8", x"78", x"0E", x"0E", x"8D", x"2D", x"0B", x"0B", x"07", x"87", x"00", x"00", x"0F", x"1F", x"1F", x"1F", x"0D", x"0D", x"00", x"00", x"0D", x"1D", x"4D", x"0D", x"52", x"32", x"05", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"9A", x"7F", x"B2", x"25", x"88", x"04", x"00", x"00", x"00", x"00", x"F0", x"F8", x"F8", x"F8", x"B8", x"B0", x"00", x"00", x"B0", x"B8", x"B8", x"B0", x"40", x"4A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04", x"04", x"08", x"08", x"FE", x"FE", x"FD", x"FD", x"FB", x"FB", x"F7", x"F7", x"10", x"10", x"20", x"20", x"40", x"40", x"80", x"80", x"EF", x"EF", x"DF", x"DF", x"BF", x"BF", x"7F", x"7F", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"C0", x"C0", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"3F", x"3F", x"00", x"00", x"00", x"00", x"FF", x"FF", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04", x"04", x"08", x"08", x"FE", x"FE", x"FD", x"FD", x"FB", x"FB", x"F7", x"F7", x"10", x"10", x"20", x"20", x"40", x"40", x"80", x"80", x"EF", x"EF", x"DF", x"DF", x"BF", x"BF", x"7F", x"7F", 
															x"DE", x"FC", x"B0", x"F0", x"E0", x"B6", x"69", x"D0", x"21", x"03", x"4F", x"0F", x"1F", x"49", x"96", x"2F", x"8C", x"80", x"80", x"00", x"81", x"80", x"8C", x"D1", x"7B", x"7F", x"7F", x"FF", x"7E", x"7F", x"73", x"2E", x"E2", x"68", x"F6", x"E0", x"B8", x"FC", x"FC", x"36", x"1D", x"97", x"09", x"1F", x"47", x"03", x"03", x"C9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5C", x"F8", x"34", x"49", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04", x"04", x"08", x"08", x"FE", x"FE", x"FD", x"FD", x"FB", x"FB", x"F7", x"F7", x"10", x"10", x"20", x"20", x"40", x"40", x"80", x"80", x"EF", x"EF", x"DF", x"DF", x"BF", x"BF", x"7F", x"7F", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"66", x"FF", x"FF", x"66", x"66", x"FF", x"FF", x"66", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"F1", x"F1", x"31", x"31", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"CF", x"CF", x"31", x"31", x"31", x"31", x"31", x"31", x"31", x"31", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"31", x"71", x"E3", x"C6", x"0C", x"18", x"F0", x"E0", x"CF", x"8F", x"1D", x"39", x"F3", x"E7", x"0F", x"1F", x"FF", x"F7", x"BF", x"00", x"EF", x"FF", x"FE", x"FF", x"00", x"08", x"40", x"FF", x"10", x"00", x"01", x"00", x"DF", x"FF", x"7D", x"FF", x"FF", x"F7", x"BF", x"00", x"20", x"00", x"82", x"00", x"00", x"08", x"40", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"4E", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"B1", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"36", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"7E", x"FF", x"FF", x"DB", x"5B", x"1A", x"00", x"00", x"7E", x"FF", x"5B", x"25", x"A4", x"E5", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"4E", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"B1", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"36", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", 
															x"38", x"9C", x"CE", x"E7", x"E7", x"CE", x"9C", x"38", x"FF", x"7F", x"3F", x"1F", x"1F", x"3F", x"7F", x"FF", x"7F", x"3F", x"1F", x"0F", x"0F", x"1F", x"3F", x"7F", x"F8", x"FC", x"FE", x"FF", x"FF", x"FE", x"FC", x"F8", x"00", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"FF", x"3F", x"1F", x"1F", x"1F", x"1F", x"1F", x"3F", x"00", x"00", x"00", x"80", x"40", x"20", x"10", x"0F", x"FF", x"FF", x"FF", x"7F", x"BF", x"DF", x"EF", x"F0", x"FE", x"01", x"01", x"01", x"01", x"01", x"01", x"FE", x"01", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"4E", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"B1", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"36", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C9", x"F3", x"CB", x"CB", x"F3", x"CB", x"CB", x"F3", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"18", x"18", x"DE", x"06", x"06", x"DC", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"06", x"38", x"C0", x"00", x"00", x"00", x"00", x"FF", x"F9", x"C7", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"1C", x"03", x"00", x"00", x"00", x"00", x"FF", x"9F", x"E3", x"FC", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"FF", x"7C", x"5C", x"5C", x"58", x"FF", x"FF", x"80", x"FF", x"7C", x"5C", x"5F", x"5F", x"58", x"5F", x"5C", x"7C", x"F8", x"80", x"80", x"FF", x"58", x"5F", x"5C", x"7C", x"FF", x"FF", x"80", x"FF", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"FE", x"FE", x"02", x"FE", x"00", x"00", x"F0", x"F0", x"10", x"F0", x"00", x"00", x"00", x"00", x"02", x"FE", x"10", x"F0", x"00", x"00", x"FE", x"FE", x"02", x"FE", x"00", x"00", x"00", x"6E", x"34", x"1E", x"0F", x"05", x"7E", x"7E", x"42", x"6E", x"34", x"1E", x"0F", x"05", x"04", x"0F", x"1E", x"3C", x"78", x"40", x"7E", x"7E", x"04", x"0F", x"1E", x"3C", x"7E", x"42", x"7E", x"7E", x"00", x"00", x"40", x"76", x"2C", x"78", x"F0", x"E0", x"7E", x"7E", x"42", x"76", x"2C", x"78", x"F0", x"E0", x"60", x"F0", x"78", x"3C", x"70", x"40", x"7E", x"7E", x"60", x"F0", x"78", x"3C", x"7E", x"42", x"7E", x"7E", 
															x"00", x"00", x"00", x"7F", x"5C", x"5C", x"5C", x"5C", x"3F", x"7F", x"40", x"7F", x"5C", x"5C", x"5C", x"5C", x"5C", x"5C", x"5C", x"5C", x"78", x"70", x"7F", x"3F", x"5C", x"5C", x"5C", x"5C", x"7F", x"70", x"7F", x"3F", x"00", x"00", x"18", x"EC", x"2E", x"3E", x"00", x"00", x"FC", x"FE", x"1E", x"EE", x"2E", x"3E", x"00", x"00", x"00", x"00", x"00", x"20", x"3E", x"1E", x"FE", x"FC", x"00", x"00", x"3E", x"3E", x"FE", x"1E", x"FE", x"FC", x"00", x"00", x"00", x"FE", x"5C", x"5C", x"5C", x"5C", x"FE", x"FE", x"82", x"FE", x"5C", x"5C", x"5C", x"5C", x"5C", x"5C", x"5C", x"5C", x"F8", x"BC", x"FE", x"FE", x"5C", x"5C", x"5C", x"5C", x"FE", x"BE", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"05", x"05", x"05", x"05", x"FF", x"FF", x"80", x"FF", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"0F", x"0B", x"0F", x"0F", x"05", x"05", x"05", x"05", x"0F", x"0B", x"0F", x"0F", 
															x"00", x"00", x"00", x"FE", x"C0", x"C0", x"C0", x"C0", x"FE", x"FE", x"02", x"FE", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"C0", x"E0", x"E0", x"C0", x"C0", x"C0", x"C0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"38", x"EC", x"2E", x"2E", x"FE", x"3C", x"FC", x"FE", x"3E", x"EE", x"2E", x"2E", x"FE", x"FC", x"3C", x"E8", x"2C", x"2E", x"EE", x"3E", x"3E", x"FC", x"3C", x"EE", x"2E", x"2E", x"EE", x"FE", x"3E", x"FC", x"80", x"00", x"BC", x"DC", x"5C", x"5C", x"5D", x"5F", x"FC", x"FC", x"BC", x"DC", x"5C", x"5C", x"5D", x"5F", x"5F", x"5D", x"5C", x"5C", x"FC", x"BC", x"FC", x"FC", x"5F", x"5D", x"5C", x"5C", x"FC", x"BC", x"FC", x"FC", x"00", x"00", x"80", x"CE", x"5C", x"F8", x"F0", x"E0", x"FE", x"FE", x"82", x"CE", x"5C", x"F8", x"F0", x"E0", x"60", x"B0", x"D8", x"5C", x"E0", x"80", x"FE", x"FE", x"60", x"B0", x"D8", x"5C", x"FE", x"86", x"FE", x"FE", 
															x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"02", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"FD", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"BF", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"02", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"FD", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"40", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"BF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", 
															x"00", x"64", x"94", x"84", x"84", x"94", x"67", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"56", x"0A", x"00", x"30", x"41", x"12", x"18", x"26", x"A9", x"F5", x"FF", x"CF", x"BE", x"FD", x"E7", x"F9", x"40", x"11", x"00", x"00", x"03", x"04", x"10", x"81", x"BF", x"EE", x"FF", x"FF", x"FC", x"FB", x"EF", x"7E", x"42", x"18", x"24", x"40", x"01", x"00", x"00", x"36", x"BD", x"E7", x"DB", x"BF", x"FE", x"FF", x"FF", x"C9", x"7F", x"3F", x"59", x"56", x"AF", x"53", x"0C", x"6B", x"80", x"C0", x"A6", x"A9", x"50", x"AC", x"F3", x"94", x"96", x"43", x"01", x"00", x"01", x"90", x"21", x"8D", x"69", x"FC", x"FE", x"FF", x"FE", x"EF", x"FE", x"72", x"53", x"07", x"6C", x"9F", x"07", x"0F", x"1F", x"76", x"AC", x"F8", x"93", x"60", x"F8", x"F0", x"E0", x"89", x"EF", x"FF", x"FE", x"FF", x"DF", x"FF", x"7D", x"FF", x"10", x"00", x"01", x"00", x"20", x"00", x"82", x"00", 
															x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"CC", x"CC", x"CC", x"CC", x"FF", x"FB", x"DF", x"FF", x"33", x"33", x"33", x"33", x"00", x"04", x"20", x"00", x"00", x"00", x"00", x"00", x"FF", x"DF", x"FD", x"FF", x"00", x"00", x"00", x"00", x"00", x"20", x"02", x"00", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"33", x"33", x"33", x"33", x"FF", x"FE", x"BF", x"FF", x"CC", x"CC", x"CC", x"CC", x"00", x"01", x"40", x"00", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"FE", x"FD", x"FB", x"F7", x"EF", x"DF", x"BF", x"7F", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", 
															x"FF", x"FF", x"FF", x"FF", x"7F", x"BF", x"DF", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"FB", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"BF", x"DF", x"EF", x"F7", x"FB", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04", x"04", x"08", x"08", x"00", x"00", x"01", x"01", x"03", x"03", x"07", x"07", x"10", x"10", x"20", x"20", x"40", x"40", x"80", x"80", x"0F", x"0F", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"01", x"01", x"02", x"02", x"04", x"04", x"08", x"08", x"FE", x"FE", x"FD", x"FD", x"FB", x"FB", x"F7", x"F7", x"10", x"10", x"20", x"20", x"40", x"40", x"80", x"80", x"EF", x"EF", x"DF", x"DF", x"BF", x"BF", x"7F", x"7F", 
															x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FD", x"FF", x"F0", x"F0", x"F4", x"F0", x"F0", x"F0", x"F2", x"F0", x"80", x"80", x"C0", x"C0", x"E0", x"E0", x"F0", x"F0", x"80", x"80", x"C0", x"C0", x"E0", x"E0", x"F0", x"F0", x"F8", x"F8", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"F8", x"F8", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"7F", x"7F", x"3F", x"3F", x"1F", x"1F", x"0F", x"0F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"07", x"03", x"03", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7E", x"3F", x"3B", x"1F", x"1F", x"0E", x"0B", x"F0", x"F1", x"F0", x"F4", x"F0", x"F0", x"F1", x"F4", x"03", x"0C", x"30", x"C0", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"03", x"0C", x"30", x"C0", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", 
															x"03", x"0C", x"30", x"C0", x"00", x"00", x"00", x"00", x"FC", x"F3", x"CF", x"3F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"03", x"0C", x"30", x"C0", x"FF", x"FF", x"FF", x"FF", x"FC", x"F3", x"CF", x"3F", x"C0", x"F0", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"C0", x"F0", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"FF", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"FF", x"3F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"0F", x"03", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", 
															x"38", x"3C", x"3C", x"3E", x"3E", x"3E", x"3F", x"3F", x"00", x"04", x"04", x"06", x"46", x"46", x"47", x"C7", x"C3", x"DF", x"DF", x"DF", x"BF", x"BF", x"BF", x"BF", x"3C", x"24", x"26", x"26", x"47", x"47", x"47", x"47", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"E0", x"E0", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"4E", x"FD", x"D8", x"FC", x"F0", x"00", x"00", x"00", x"B1", x"02", x"27", x"03", x"0F", 
															x"FF", x"FF", x"FF", x"4E", x"CB", x"80", x"28", x"00", x"00", x"00", x"00", x"B1", x"34", x"7F", x"DF", x"FF", x"FF", x"FF", x"FF", x"4E", x"BF", x"9F", x"0D", x"27", x"00", x"00", x"00", x"B1", x"40", x"E0", x"F2", x"D8", x"F0", x"F8", x"D2", x"6E", x"FF", x"FF", x"FF", x"FF", x"0F", x"07", x"2D", x"91", x"00", x"00", x"00", x"00", x"02", x"80", x"10", x"B5", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"EF", x"4A", x"00", x"00", x"00", x"00", x"17", x"83", x"0E", x"DC", x"FF", x"FF", x"FF", x"FF", x"E8", x"7C", x"F1", x"23", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"1C", x"38", x"70", x"E0", x"00", x"00", x"04", x"0C", x"1C", x"38", x"70", x"E0", x"00", x"00", x"E0", x"70", x"38", x"1C", x"0F", x"07", x"03", x"00", x"E0", x"70", x"38", x"1C", x"0F", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", 
															x"00", x"40", x"60", x"70", x"38", x"1C", x"0E", x"00", x"00", x"40", x"60", x"70", x"38", x"1C", x"0E", x"00", x"00", x"0E", x"1C", x"38", x"70", x"E0", x"C0", x"80", x"00", x"0E", x"1C", x"38", x"70", x"E0", x"C0", x"80", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"04", x"04", x"EE", x"84", x"64", x"24", x"E4", x"00", x"04", x"04", x"EE", x"84", x"64", x"24", x"E4", x"00", x"02", x"02", x"EE", x"AA", x"AA", x"AA", x"AE", x"00", x"02", x"02", x"EE", x"AA", x"AA", x"AA", x"AE", x"00", x"02", x"02", x"EE", x"AA", x"8A", x"8A", x"8E", x"00", x"02", x"02", x"EE", x"AA", x"8A", x"8A", x"8E", x"00", x"48", x"48", x"EE", x"4A", x"4A", x"4A", x"4A", x"00", x"48", x"48", x"EE", x"4A", x"4A", x"4A", x"4A", x"00", x"48", x"48", x"EE", x"4A", x"4A", x"4A", x"4A", x"00", x"48", x"48", x"EE", x"4A", x"4A", x"4A", x"4A", x"00", 
															x"00", x"7C", x"00", x"00", x"00", x"7C", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"18", x"08", x"10", x"20", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0C", x"1C", x"1C", x"18", x"10", x"00", x"20", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"18", x"18", x"00", x"00", x"18", x"18", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF");
	
	constant MS_PAC_MAN_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"01", x"1F", x"1F", x"0E", x"0D", x"3F", x"0C", x"0E", x"0E", x"18", x"78", x"70", x"31", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"70", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"00", x"00", x"3C", x"3F", x"3B", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"F8", x"E0", x"00", x"00", x"00", x"00", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"1F", x"1E", x"0D", x"0D", x"3E", x"0C", x"0E", x"0E", x"18", x"78", x"71", x"30", x"00", x"00", x"00", x"E0", x"C0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"3C", x"3E", x"3B", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"00", 
															x"00", x"00", x"01", x"1F", x"1F", x"0F", x"08", x"3F", x"0C", x"0E", x"0E", x"18", x"78", x"70", x"30", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FC", x"7E", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"3F", x"3F", x"3B", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"FC", x"FE", x"FC", x"FC", x"F8", x"E0", x"00", x"06", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"01", x"E7", x"0F", x"8E", x"0D", x"3F", x"0C", x"0E", x"0E", x"18", x"70", x"70", x"31", x"00", x"00", x"F0", x"01", x"E7", x"0E", x"8D", x"0D", x"3E", x"0C", x"0E", x"0E", x"18", x"70", x"71", x"30", x"00", x"00", x"F0", x"01", x"E7", x"0F", x"8F", x"08", x"3F", x"0C", x"0E", x"0E", x"18", x"70", x"70", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"07", x"1F", x"3F", x"3B", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"98", x"F8", x"F8", x"B8", x"DC", x"00", x"30", x"70", x"78", x"1F", x"07", x"06", x"40", x"7C", x"7C", x"78", x"38", x"30", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"5C", x"7C", x"3C", x"38", x"18", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"00", x"00", x"00", x"00", x"07", x"1F", x"3F", x"3B", x"7E", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"98", x"F8", x"F8", x"98", x"6C", x"00", x"30", x"70", x"78", x"1F", x"07", x"06", x"20", x"78", x"70", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"3C", x"1C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"07", x"1F", x"3F", x"3B", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"98", x"F8", x"B8", x"B8", x"BC", x"00", x"30", x"70", x"78", x"1F", x"07", x"06", x"00", x"7F", x"7F", x"7F", x"3F", x"3F", x"1E", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"BC", x"FC", x"FC", x"F8", x"F8", x"F0", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"2A", x"0A", x"8A", x"82", x"F0", x"F8", x"B8", x"DC", x"00", x"30", x"70", x"78", x"0F", x"07", x"06", x"40", x"2A", x"0A", x"8A", x"82", x"F0", x"F8", x"98", x"6C", x"00", x"30", x"70", x"78", x"0F", x"07", x"06", x"20", x"2A", x"0A", x"8A", x"82", x"F0", x"F8", x"B8", x"BC", x"00", x"30", x"70", x"78", x"0F", x"07", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"03", x"03", x"13", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"0C", x"1E", x"1E", x"1E", x"0C", x"00", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"00", x"00", x"00", x"0C", x"1E", x"1E", x"73", x"73", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"1E", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"0F", x"4F", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"3C", x"00", x"C0", x"F0", x"F8", x"FC", x"FC", x"3C", x"3E", x"00", x"00", x"00", x"00", x"60", x"F0", x"F0", x"F0", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"76", x"62", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"73", x"73", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"1E", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"DE", x"8C", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"00", x"19", x"26", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"00", x"19", x"26", x"00", x"00", x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FD", x"FD", x"FD", x"81", x"FF", x"00", x"06", x"06", x"06", x"06", x"7E", x"7E", x"00", 
															x"00", x"00", x"0C", x"1E", x"1E", x"1E", x"0C", x"00", x"00", x"03", x"03", x"13", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"1E", x"1E", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"1E", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"73", x"73", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"3C", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"0F", x"4F", x"00", x"00", x"00", x"00", x"60", x"F0", x"F0", x"F0", x"00", x"C0", x"F0", x"F8", x"FC", x"FC", x"3C", x"3E", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"76", x"62", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"1E", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"73", x"73", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"DE", x"8C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"00", x"19", x"26", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"00", x"19", x"26", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"00", x"12", x"1E", x"1E", x"0C", x"00", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"12", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"00", x"00", x"00", x"00", x"18", x"3C", x"0C", x"0C", x"00", x"C0", x"F0", x"F8", x"FC", x"FC", x"FC", x"FE", x"00", x"00", x"00", x"00", x"60", x"F0", x"30", x"30", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"12", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"3F", x"7F", x"00", x"03", x"0F", x"1F", x"3F", x"39", x"39", x"7F", x"7F", x"7F", x"7F", x"7F", x"6E", x"46", x"00", x"00", x"7F", x"66", x"59", x"7F", x"6E", x"46", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7B", x"31", x"00", x"00", x"7F", x"66", x"59", x"7F", x"7B", x"31", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"20", x"20", x"EE", x"2A", x"2A", x"EA", x"0A", x"E0", x"20", x"20", x"EE", x"2A", x"2A", x"EA", x"0A", x"80", x"A0", x"A0", x"EE", x"2A", x"2A", x"2A", x"0A", x"80", x"A0", x"A0", x"EE", x"2A", x"2A", x"2A", x"0A", x"E0", x"A0", x"A0", x"EE", x"AA", x"AA", x"EA", x"0A", x"E0", x"A0", x"A0", x"EE", x"AA", x"AA", x"EA", x"0A", x"E0", x"A0", x"A0", x"EE", x"2A", x"2A", x"2A", x"0A", x"E0", x"A0", x"A0", x"EE", x"2A", x"2A", x"2A", x"0A", 
															x"E0", x"80", x"80", x"EE", x"2A", x"2A", x"EA", x"0A", x"E0", x"80", x"80", x"EE", x"2A", x"2A", x"EA", x"0A", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"A0", x"0A", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"0A", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"A0", x"AE", x"AA", x"AA", x"EA", x"0A", x"0A", x"0E", x"A0", x"AE", x"AA", x"AA", x"EA", x"0A", x"0A", x"0E", x"E0", x"20", x"20", x"EE", x"8A", x"8A", x"EA", x"0A", x"E0", x"20", x"20", x"EE", x"8A", x"8A", x"EA", x"0A", x"40", x"40", x"40", x"4E", x"4A", x"4A", x"4A", x"0A", x"40", x"40", x"40", x"4E", x"4A", x"4A", x"4A", x"0A", x"00", x"00", x"00", x"0E", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"0E", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"0E", x"08", x"08", x"0E", x"02", x"00", x"00", x"00", x"0E", x"08", x"08", x"0E", x"02", x"02", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"02", x"02", x"0E", x"08", x"00", x"00", x"00", x"0E", x"02", x"02", x"0E", x"08", x"08", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"04", x"04", x"04", x"00", x"00", x"00", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"EE", x"AA", x"AA", x"EA", x"0A", x"80", x"80", x"80", x"EE", x"AA", x"AA", x"EA", x"0A", x"E0", x"20", x"20", x"2E", x"2A", x"2A", x"2A", x"0A", x"E0", x"20", x"20", x"2E", x"2A", x"2A", x"2A", x"0A", 
															x"18", x"25", x"25", x"05", x"09", x"11", x"21", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"29", x"29", x"29", x"29", x"29", x"29", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"19", x"29", x"49", x"7D", x"09", x"09", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"25", x"25", x"19", x"25", x"25", x"25", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"98", x"A5", x"A1", x"B9", x"A5", x"A5", x"A5", x"98", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"18", x"3C", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"24", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"60", x"F0", x"F0", x"F0", x"60", x"00", x"00", x"00", x"60", x"F0", x"30", x"30", x"60", x"00", x"00", x"00", x"24", x"3C", x"3C", x"18", x"00", x"00", x"00", x"18", x"3C", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"60", x"F0", x"30", x"30", x"60", x"00", x"00", x"00", x"60", x"F0", x"F0", x"F0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"25", x"25", x"05", x"09", x"11", x"21", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"29", x"29", x"29", x"29", x"29", x"29", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"19", x"29", x"49", x"7D", x"09", x"09", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"25", x"25", x"19", x"25", x"25", x"25", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"98", x"A5", x"A1", x"B9", x"A5", x"A5", x"A5", x"98", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"77", x"24", x"26", x"24", x"27", x"00", x"00", x"00", x"77", x"24", x"26", x"24", x"27", x"00", x"00", x"00", x"4B", x"6B", x"5B", x"48", x"4B", x"00", x"00", x"00", x"4B", x"6B", x"5B", x"48", x"4B", x"00", x"00", x"31", x"4A", x"4A", x"4A", x"4A", x"4A", x"31", x"00", x"31", x"4A", x"4A", x"4A", x"4A", x"4A", x"31", x"00", x"8C", x"52", x"52", x"52", x"52", x"52", x"8C", x"00", x"8C", x"52", x"52", x"52", x"52", x"52", x"8C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"1C", x"3A", x"3E", x"3D", x"00", x"00", x"00", x"01", x"02", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B0", x"B8", x"00", x"18", x"78", x"90", x"10", x"20", x"40", x"40", x"3D", x"3D", x"3D", x"1D", x"01", x"00", x"00", x"00", x"00", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"B8", x"B8", x"F8", x"F8", x"F8", x"F0", x"00", x"00", x"40", x"40", x"00", x"80", x"40", x"00", x"00", x"00", x"00", x"01", x"00", x"18", x"3C", x"3F", x"3F", x"3F", x"00", x"01", x"0F", x"07", x"03", x"10", x"05", x"00", x"00", x"00", x"10", x"38", x"78", x"F8", x"F8", x"F8", x"00", x"00", x"E0", x"C0", x"90", x"40", x"00", x"20", x"1F", x"1F", x"1F", x"07", x"01", x"00", x"00", x"00", x"01", x"08", x"02", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"1C", x"3E", x"3E", x"7F", x"7F", x"7F", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"38", x"FC", x"FE", x"FE", x"FE", x"FE", x"80", x"80", x"00", x"10", x"00", x"00", x"00", x"10", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"3E", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"F8", x"70", x"10", x"30", x"20", x"60", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"0F", x"1F", x"3F", x"3F", x"00", x"60", x"F8", x"F8", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"F8", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"1F", x"1F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"F8", x"F8", x"E0", x"00", x"00", x"00", 
															x"00", x"60", x"00", x"00", x"00", x"00", x"20", x"10", x"18", x"7C", x"76", x"66", x"60", x"61", x"61", x"73", x"00", x"00", x"84", x"00", x"00", x"00", x"01", x"22", x"1C", x"3E", x"E6", x"C3", x"C3", x"83", x"83", x"23", x"00", x"00", x"00", x"00", x"00", x"20", x"30", x"00", x"32", x"16", x"04", x"1C", x"19", x"71", x"F0", x"40", x"00", x"00", x"00", x"00", x"00", x"06", x"00", x"00", x"67", x"76", x"34", x"10", x"D8", x"CE", x"06", x"00", x"00", x"00", x"00", x"02", x"07", x"07", x"07", x"0F", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"0F", x"07", x"00", x"00", x"00", x"04", x"04", x"02", x"00", x"00", x"E0", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"30", x"38", x"38", x"78", x"F8", x"F0", x"00", x"00", x"10", x"20", x"00", x"00", x"40", x"80", x"03", x"07", x"0F", x"1F", x"3F", x"FE", x"78", x"00", x"01", x"02", x"04", x"08", x"10", x"00", x"00", x"00", x"F0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"08", x"10", x"20", x"20", x"20", x"00", x"07", x"1F", x"3C", x"30", x"70", x"60", x"60", x"0E", x"1F", x"1F", x"6F", x"F7", x"FE", x"FC", x"79", x"0E", x"1F", x"1F", x"6F", x"F4", x"F9", x"F3", x"76", x"3F", x"3F", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"0C", x"07", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"E0", x"00", x"00", x"18", x"F0", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3F", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"F8", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3E", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FC", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FC", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"3E", x"3C", x"1C", x"18", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"3E", x"1E", x"1C", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FC", x"7E", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"38", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"0E", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FC", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"3F", x"3F", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"07", x"0C", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"E0", x"00", x"00", x"00", x"F0", x"18", x"00", x"00", x"00", x"00", 
															x"00", x"FC", x"03", x"EF", x"1F", x"DF", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"15", x"15", x"E5", x"F9", x"FD", x"FD", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"15", x"15", x"E5", x"F9", x"FD", x"FD", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"F8", x"E0", x"E0", x"F8", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"34", x"39", x"06", x"1F", x"1F", x"3F", x"3F", x"19", x"2B", x"3E", x"19", x"00", x"03", x"03", x"00", x"00", x"40", x"0C", x"30", x"FC", x"FC", x"FE", x"FE", x"CC", x"BE", x"FE", x"CC", x"00", x"60", x"60", x"00", x"00", x"42", x"C3", x"E7", x"E7", x"FF", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"E7", x"E7", x"C3", x"42", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"C0", x"F8", x"C0", x"C0", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"6C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"CC", x"CC", x"CC", x"78", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"38", x"30", x"20", x"00", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"36", x"62", x"43", x"C0", x"80", x"80", x"80", x"1C", x"3E", x"7E", x"7F", x"FF", x"FF", x"FF", x"FF", x"C0", x"40", x"60", x"20", x"30", x"1C", x"06", x"03", x"FF", x"7F", x"7F", x"3F", x"3F", x"1F", x"07", x"03", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"FE", x"FE", x"FE", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"74", x"FF", x"FF", x"3F", x"00", x"00", x"00", x"1C", x"7C", x"FF", x"FF", x"3F", x"00", x"00", x"03", x"0F", x"3F", x"7F", x"FF", x"FF", x"FF", x"00", x"03", x"0F", x"3F", x"7F", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"01", x"06", x"1F", x"11", x"3F", x"00", x"00", x"00", x"01", x"06", x"1F", x"11", x"3F", x"01", x"06", x"1F", x"61", x"FE", x"18", x"E0", x"80", x"01", x"06", x"1F", x"61", x"FE", x"18", x"E0", x"80", x"00", x"06", x"1F", x"61", x"FE", x"18", x"E0", x"80", x"00", x"06", x"1F", x"61", x"FE", x"18", x"E0", x"80", x"00", x"00", x"00", x"07", x"3C", x"3F", x"38", x"3F", x"00", x"00", x"00", x"07", x"3C", x"3F", x"38", x"3F", x"03", x"1F", x"F0", x"FF", x"07", x"FC", x"E0", x"00", x"03", x"1F", x"F0", x"FF", x"07", x"FC", x"E0", x"00", x"01", x"0F", x"7F", x"C0", x"FF", x"1E", x"F0", x"80", x"01", x"0F", x"7F", x"C0", x"FF", x"1E", x"F0", x"80", x"00", x"06", x"3A", x"FF", x"03", x"FF", x"78", x"C0", x"00", x"06", x"3A", x"FF", x"03", x"FF", x"78", x"C0", x"00", x"00", x"00", x"00", x"3F", x"26", x"33", x"39", x"00", x"00", x"00", x"00", x"3F", x"26", x"33", x"39", 
															x"00", x"00", x"00", x"00", x"FF", x"66", x"33", x"99", x"00", x"00", x"00", x"00", x"FF", x"66", x"33", x"99", x"00", x"00", x"00", x"00", x"C0", x"40", x"40", x"C0", x"00", x"00", x"00", x"00", x"C0", x"40", x"40", x"C0", x"FC", x"F8", x"F0", x"E0", x"C0", x"C0", x"E0", x"FC", x"FC", x"F8", x"F0", x"E0", x"C0", x"C0", x"E0", x"FC", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FE", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"FE", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"80", x"E0", x"FC", x"00", x"00", x"00", x"00", x"00", x"80", x"E0", x"FC", x"FF", x"FF", x"FF", x"7F", x"7F", x"3E", x"1C", x"08", x"FF", x"FF", x"FF", x"7F", x"7F", x"3E", x"1C", x"08", 
															x"00", x"00", x"00", x"07", x"0F", x"1F", x"3F", x"3F", x"70", x"78", x"7F", x"78", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FE", x"FE", x"07", x"1F", x"FF", x"1F", x"07", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"C3", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"7C", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"38", x"7C", x"7C", x"38", x"00", x"00", x"00", x"44", x"44", x"00", x"00", x"00", x"00", x"00", x"99", x"5A", x"00", x"C3", x"C3", x"00", x"5A", x"99", x"99", x"5A", x"00", x"C3", x"C3", x"00", x"5A", x"99", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", 
															x"38", x"7C", x"FE", x"FE", x"BE", x"3E", x"1C", x"00", x"38", x"7C", x"FE", x"FE", x"BE", x"3E", x"1C", x"00", x"07", x"0F", x"1F", x"1F", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"00", x"00", x"07", x"07", x"03", x"03", x"01", x"01", x"1F", x"0F", x"07", x"07", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"0F", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"10", x"10", x"30", x"30", x"30", x"60", x"60", x"00", x"C0", x"C0", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"71", x"73", x"36", x"3C", x"E9", x"F2", x"7C", x"7F", x"51", x"52", x"55", x"5A", x"94", x"89", x"82", x"80", x"80", x"60", x"40", x"B0", x"20", x"50", x"A0", x"40", x"00", x"C0", x"20", x"70", x"90", x"30", x"60", x"C0", x"7E", x"7D", x"7D", x"3C", x"9F", x"81", x"8E", x"4C", x"81", x"83", x"83", x"C3", x"E0", x"FE", x"FF", x"7C", x"80", x"00", x"00", x"80", x"00", x"80", x"80", x"00", x"80", x"00", x"00", x"80", x"80", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"30", x"18", x"00", x"00", x"00", x"00", x"70", x"F8", x"FC", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"37", x"33", x"31", x"30", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"0F", x"07", x"03", x"01", x"07", x"0C", x"18", x"10", x"10", x"18", x"0C", x"07", x"07", x"0C", x"18", x"10", x"10", x"18", x"0C", x"07", x"01", x"03", x"03", x"07", x"0F", x"FF", x"FF", x"7F", x"00", x"01", x"01", x"03", x"03", x"07", x"79", x"3A", x"E0", x"F0", x"F0", x"F8", x"F8", x"FF", x"FF", x"FF", x"00", x"80", x"80", x"C0", x"C0", x"E0", x"BE", x"5C", x"3F", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"7C", x"19", x"0B", x"0B", x"1F", x"1E", x"38", x"20", x"00", x"FF", x"FE", x"FC", x"FE", x"FE", x"FF", x"1F", x"07", x"18", x"50", x"50", x"F8", x"78", x"1C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"3C", x"7E", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E3", x"C1", x"83", x"8F", x"8F", x"83", x"C1", x"E3", x"1C", x"3E", x"7C", x"70", x"70", x"7C", x"3E", x"1C", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"81", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"81", x"FF", x"00", x"FF", x"81", x"BD", x"BD", x"BD", x"BD", x"81", x"FF", x"00", x"7E", x"7E", x"66", x"66", x"7E", x"7E", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"1C", x"3A", x"3E", x"3D", x"00", x"00", x"00", x"01", x"02", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B0", x"B8", x"00", x"18", x"78", x"90", x"10", x"20", x"40", x"40", x"3D", x"3D", x"3D", x"1D", x"01", x"00", x"00", x"00", x"00", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"B8", x"B8", x"F8", x"F8", x"F8", x"F0", x"00", x"00", x"40", x"40", x"00", x"80", x"40", x"00", x"00", x"00", x"00", x"01", x"00", x"18", x"3C", x"3F", x"3F", x"3F", x"00", x"01", x"0F", x"07", x"03", x"10", x"05", x"00", x"00", x"00", x"10", x"38", x"78", x"F8", x"F8", x"F8", x"00", x"00", x"E0", x"C0", x"90", x"40", x"00", x"20", x"1F", x"1F", x"1F", x"07", x"01", x"00", x"00", x"00", x"01", x"08", x"02", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"1C", x"3E", x"3E", x"7F", x"7F", x"7F", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"38", x"FC", x"FE", x"FE", x"FE", x"FE", x"80", x"80", x"00", x"10", x"00", x"00", x"00", x"10", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"3E", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"F8", x"70", x"10", x"30", x"20", x"60", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"0F", x"1F", x"3F", x"3F", x"00", x"60", x"F8", x"F8", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"F8", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"1F", x"1F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"F8", x"F8", x"E0", x"00", x"00", x"00", 
															x"00", x"60", x"00", x"00", x"00", x"00", x"20", x"10", x"18", x"7C", x"76", x"66", x"60", x"61", x"61", x"73", x"00", x"00", x"84", x"00", x"00", x"00", x"01", x"22", x"1C", x"3E", x"E6", x"C3", x"C3", x"83", x"83", x"23", x"00", x"00", x"00", x"00", x"00", x"20", x"30", x"00", x"32", x"16", x"04", x"1C", x"19", x"71", x"F0", x"40", x"00", x"00", x"00", x"00", x"00", x"06", x"00", x"00", x"67", x"76", x"34", x"10", x"D8", x"CE", x"06", x"00", x"00", x"00", x"00", x"02", x"07", x"07", x"07", x"0F", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"0F", x"07", x"00", x"00", x"00", x"04", x"04", x"02", x"00", x"00", x"E0", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"30", x"38", x"38", x"78", x"F8", x"F0", x"00", x"00", x"10", x"20", x"00", x"00", x"40", x"80", x"03", x"07", x"0F", x"1F", x"3F", x"FE", x"78", x"00", x"01", x"02", x"04", x"08", x"10", x"00", x"00", x"00", x"F0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"0F", x"0F", x"0F", x"3F", x"0C", x"0E", x"0E", x"18", x"71", x"73", x"32", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"F0", x"C0", x"00", x"00", x"00", x"00", x"04", x"80", x"00", x"00", x"00", x"3C", x"3F", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"F8", x"E0", x"00", x"00", x"00", x"00", x"0C", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"07", x"1F", x"3F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"F8", x"F8", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", x"1F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FC", x"FC", x"F8", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"70", x"60", x"60", x"60", x"70", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"0E", x"06", x"06", x"06", x"0E", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"7C", x"00", x"3C", x"00", x"1C", x"00", x"00", x"FF", x"7C", x"00", x"3C", x"00", x"1C", x"FF", x"00", x"00", x"8A", x"DA", x"AA", x"8A", x"8A", x"00", x"00", x"FF", x"8A", x"DA", x"AA", x"8A", x"8A", x"FF", x"00", x"00", x"8A", x"CA", x"AA", x"9A", x"8A", x"00", x"00", x"FF", x"8A", x"CA", x"AA", x"9A", x"8A", x"FF", x"00", x"00", x"39", x"25", x"39", x"25", x"39", x"00", x"00", x"FF", x"39", x"25", x"39", x"25", x"39", x"FF", x"00", x"00", x"3C", x"20", x"2C", x"24", x"3C", x"00", x"00", x"FF", x"3C", x"20", x"2C", x"24", x"3C", x"FF", x"00", x"00", x"FF", x"8A", x"EB", x"2A", x"EA", x"00", x"00", x"FF", x"FF", x"8A", x"EB", x"2A", x"EA", x"FF", x"00", x"00", x"39", x"AD", x"3B", x"A9", x"A9", x"00", x"00", x"FF", x"39", x"AD", x"3B", x"A9", x"A9", x"FF", x"00", x"00", x"77", x"44", x"56", x"54", x"77", x"00", x"00", x"FF", x"77", x"44", x"56", x"54", x"77", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"07", x"00", x"00", x"00", x"00", x"03", x"04", x"08", x"08", x"07", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"03", x"00", x"00", x"00", x"00", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"FF", x"FF", x"FF", x"F8", x"F0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"07", x"08", x"10", x"10", x"10", x"07", x"07", x"07", x"0F", x"1F", x"FF", x"FF", x"FF", x"08", x"08", x"08", x"10", x"E0", x"00", x"00", x"00", x"00", x"0F", x"3F", x"38", x"70", x"60", x"60", x"60", x"0F", x"30", x"40", x"47", x"88", x"90", x"90", x"90", x"60", x"60", x"60", x"70", x"38", x"3F", x"0F", x"00", x"90", x"90", x"90", x"88", x"47", x"40", x"30", x"0F", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"90", x"90", x"90", x"90", x"90", x"90", x"90", x"90", 
															x"00", x"FF", x"FF", x"F8", x"F0", x"E0", x"E0", x"E0", x"FF", x"00", x"00", x"07", x"08", x"10", x"10", x"10", x"7F", x"7F", x"7F", x"78", x"70", x"60", x"60", x"60", x"80", x"80", x"80", x"87", x"88", x"90", x"90", x"90", x"07", x"07", x"07", x"0F", x"1F", x"FF", x"FF", x"00", x"08", x"08", x"08", x"10", x"E0", x"00", x"00", x"FF", x"06", x"06", x"06", x"0E", x"1E", x"FE", x"FE", x"FE", x"09", x"09", x"09", x"11", x"E1", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"06", x"00", x"00", x"00", x"00", x"0F", x"08", x"08", x"09", x"06", x"07", x"07", x"00", x"00", x"00", x"00", x"00", x"09", x"08", x"08", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"FF", x"01", x"01", x"FF", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"FF", x"80", x"80", x"80", 
															x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"06", x"06", x"00", x"00", x"00", x"00", x"03", x"05", x"09", x"09", x"06", x"06", x"02", x"00", x"00", x"00", x"00", x"00", x"09", x"09", x"05", x"03", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"0E", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0E", x"FF", x"8B", x"AB", x"8B", x"BB", x"BB", x"B8", x"FF", x"00", x"74", x"54", x"74", x"44", x"44", x"47", x"00", x"FF", x"8A", x"AA", x"88", x"AD", x"AD", x"AD", x"FF", x"00", x"75", x"55", x"77", x"52", x"52", x"52", x"00", x"FF", x"D1", x"D5", x"CD", x"CD", x"D5", x"D4", x"FF", x"00", x"2E", x"2A", x"32", x"32", x"2A", x"2B", x"00", x"FF", x"82", x"AA", x"8D", x"AD", x"AA", x"2A", x"FF", x"00", x"7D", x"55", x"72", x"52", x"55", x"D5", x"00", 
															x"00", x"00", x"00", x"00", x"03", x"07", x"0C", x"0D", x"00", x"00", x"00", x"00", x"03", x"04", x"0B", x"0B", x"0D", x"0C", x"07", x"03", x"00", x"00", x"00", x"00", x"0B", x"0B", x"04", x"03", x"00", x"00", x"00", x"00", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"FF", x"80", x"9F", x"BF", x"B8", x"B0", x"B0", x"B0", x"FF", x"FF", x"E0", x"CF", x"D8", x"D0", x"D0", x"D0", x"0D", x"0D", x"0D", x"1D", x"FD", x"F9", x"01", x"FF", x"0B", x"0B", x"0B", x"1B", x"F3", x"07", x"FF", x"FF", x"FF", x"03", x"03", x"CF", x"CC", x"CD", x"CC", x"FF", x"00", x"FC", x"FC", x"30", x"33", x"32", x"33", x"00", x"FF", x"FD", x"FD", x"FD", x"44", x"55", x"44", x"FF", x"00", x"02", x"02", x"02", x"BB", x"AA", x"BB", x"00", x"FF", x"FC", x"FE", x"FF", x"51", x"55", x"55", x"FF", x"00", x"03", x"01", x"00", x"AE", x"AA", x"AA", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"C0", x"20", x"10", x"10", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"20", x"C0", x"00", x"00", x"00", x"00", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"FF", x"FF", x"1F", x"0F", x"07", x"07", x"07", x"00", x"00", x"00", x"E0", x"10", x"08", x"08", x"08", x"E0", x"E0", x"E0", x"F0", x"F8", x"FF", x"FF", x"FF", x"10", x"10", x"10", x"08", x"07", x"00", x"00", x"00", x"00", x"F0", x"FC", x"1C", x"0E", x"06", x"06", x"06", x"F0", x"0C", x"02", x"E2", x"11", x"09", x"09", x"09", x"06", x"06", x"06", x"0E", x"1C", x"FC", x"F0", x"00", x"09", x"09", x"09", x"11", x"E2", x"02", x"0C", x"F0", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", 
															x"00", x"FF", x"FF", x"1F", x"0F", x"07", x"07", x"07", x"FF", x"00", x"00", x"E0", x"10", x"08", x"08", x"08", x"FE", x"FE", x"FE", x"1E", x"0E", x"06", x"06", x"06", x"01", x"01", x"01", x"E1", x"11", x"09", x"09", x"09", x"E0", x"E0", x"E0", x"F0", x"F8", x"FF", x"FF", x"00", x"10", x"10", x"10", x"08", x"07", x"00", x"00", x"FF", x"60", x"60", x"60", x"70", x"78", x"7F", x"7F", x"7F", x"90", x"90", x"90", x"88", x"87", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"60", x"00", x"00", x"00", x"00", x"F0", x"10", x"10", x"90", x"60", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"90", x"10", x"10", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"FF", x"80", x"80", x"FF", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"FF", x"01", x"01", x"01", 
															x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"60", x"60", x"00", x"00", x"00", x"00", x"C0", x"A0", x"90", x"90", x"60", x"60", x"40", x"00", x"00", x"00", x"00", x"00", x"90", x"90", x"A0", x"C0", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"70", x"50", x"50", x"50", x"50", x"50", x"50", x"70", x"FF", x"82", x"AA", x"8D", x"AD", x"AA", x"2A", x"FF", x"00", x"7D", x"55", x"72", x"52", x"55", x"D5", x"00", x"FF", x"D1", x"D5", x"CD", x"CD", x"D5", x"D4", x"FF", x"00", x"2E", x"2A", x"32", x"32", x"2A", x"2B", x"00", x"FF", x"8A", x"AA", x"88", x"AD", x"AD", x"AD", x"FF", x"00", x"75", x"55", x"77", x"52", x"52", x"52", x"00", x"FF", x"8B", x"AB", x"8B", x"BB", x"BB", x"B8", x"FF", x"00", x"74", x"54", x"74", x"44", x"44", x"47", x"00", 
															x"00", x"00", x"00", x"00", x"C0", x"E0", x"30", x"B0", x"00", x"00", x"00", x"00", x"C0", x"20", x"D0", x"D0", x"B0", x"30", x"E0", x"C0", x"00", x"00", x"00", x"00", x"D0", x"D0", x"20", x"C0", x"00", x"00", x"00", x"00", x"B0", x"B0", x"B0", x"B0", x"B0", x"B0", x"B0", x"B0", x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"D0", x"FF", x"01", x"F9", x"FD", x"1D", x"0D", x"0D", x"0D", x"FF", x"FF", x"07", x"F3", x"1B", x"0B", x"0B", x"0B", x"B0", x"B0", x"B0", x"B8", x"BF", x"9F", x"80", x"FF", x"D0", x"D0", x"D0", x"D8", x"CF", x"E0", x"FF", x"FF", x"FF", x"FC", x"FE", x"FF", x"51", x"55", x"55", x"FF", x"00", x"03", x"01", x"00", x"AE", x"AA", x"AA", x"00", x"FF", x"FD", x"FD", x"FD", x"44", x"55", x"44", x"FF", x"00", x"02", x"02", x"02", x"BB", x"AA", x"BB", x"00", x"FF", x"03", x"03", x"CF", x"CC", x"CD", x"CC", x"FF", x"00", x"FC", x"FC", x"30", x"33", x"32", x"33", x"00", 
															x"00", x"38", x"44", x"C6", x"C6", x"C6", x"44", x"38", x"00", x"38", x"44", x"C6", x"C6", x"C6", x"44", x"38", x"00", x"30", x"70", x"30", x"30", x"30", x"30", x"FC", x"00", x"30", x"70", x"30", x"30", x"30", x"30", x"FC", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"FE", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"FE", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", 
															x"00", x"78", x"C4", x"E4", x"78", x"9E", x"86", x"7C", x"00", x"78", x"C4", x"E4", x"78", x"9E", x"86", x"7C", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00", x"30", x"30", x"10", x"20", x"00", x"00", x"00", x"00", x"30", x"30", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"10", x"20", x"40", x"20", x"10", x"00", x"00", x"00", x"10", x"20", x"40", x"20", x"10", x"00", x"00", x"1C", x"3C", x"38", x"30", x"20", x"00", x"40", x"00", x"1C", x"3C", x"38", x"30", x"20", x"00", x"40", x"18", x"0C", x"06", x"FF", x"FF", x"06", x"0C", x"18", x"18", x"0C", x"06", x"FF", x"FF", x"06", x"0C", x"18", x"00", x"7C", x"C6", x"0C", x"18", x"00", x"18", x"18", x"00", x"7C", x"C6", x"0C", x"18", x"00", x"18", x"18", 
															x"00", x"38", x"44", x"BA", x"A2", x"BA", x"44", x"38", x"00", x"38", x"44", x"BA", x"A2", x"BA", x"44", x"38", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"FC", x"C0", x"C0", x"F8", x"C0", x"C0", x"FC", x"00", x"FC", x"C0", x"C0", x"F8", x"C0", x"C0", x"FC", x"00", x"FC", x"C0", x"C0", x"F8", x"C0", x"C0", x"C0", x"00", x"FC", x"C0", x"C0", x"F8", x"C0", x"C0", x"C0", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", 
															x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"FC", x"30", x"30", x"30", x"30", x"30", x"FC", x"00", x"FC", x"30", x"30", x"30", x"30", x"30", x"FC", x"00", x"06", x"06", x"06", x"06", x"06", x"C6", x"7C", x"00", x"06", x"06", x"06", x"06", x"06", x"C6", x"7C", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FC", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FC", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", 
															x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"7C", x"C6", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"7C", x"C6", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"FC", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"FC", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"C6", x"C6", x"C6", x"EE", x"6C", x"38", x"10", x"00", x"C6", x"C6", x"C6", x"EE", x"6C", x"38", x"10", x"00", x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", 
															x"00", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"CC", x"CC", x"CC", x"78", x"30", x"30", x"30", x"00", x"CC", x"CC", x"CC", x"78", x"30", x"30", x"30", x"00", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"D8", x"D8", x"90", x"48", x"00", x"00", x"00", x"00", x"D8", x"D8", x"90", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"38", x"00", x"00", x"00", x"00", x"36", x"36", x"12", x"24", x"00", x"00", x"00", x"00", x"36", x"36", x"12", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FD", x"FD", x"FD", x"81", x"FF", x"00", x"02", x"02", x"02", x"02", x"02", x"7E", x"00", 
															x"00", x"00", x"3F", x"19", x"0B", x"0E", x"0F", x"08", x"00", x"00", x"3F", x"19", x"0B", x"0E", x"0F", x"08", x"00", x"00", x"FF", x"99", x"33", x"66", x"FF", x"00", x"00", x"00", x"FF", x"99", x"33", x"66", x"FF", x"00", x"00", x"00", x"C0", x"C0", x"40", x"40", x"C0", x"40", x"00", x"00", x"C0", x"C0", x"40", x"40", x"C0", x"40", x"08", x"09", x"09", x"0B", x"0B", x"0A", x"0A", x"0A", x"08", x"09", x"09", x"0B", x"0B", x"0A", x"0A", x"0A", x"87", x"CC", x"48", x"68", x"E8", x"28", x"2C", x"27", x"87", x"CC", x"48", x"68", x"E8", x"28", x"2C", x"27", x"7C", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"7C", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"08", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AE", x"AA", x"EE", x"AA", x"AA", x"00", x"00", x"FF", x"AE", x"AA", x"EE", x"AA", x"AA", x"FF", x"00", x"00", x"CC", x"AA", x"CA", x"AA", x"AC", x"00", x"00", x"FF", x"CC", x"AA", x"CA", x"AA", x"AC", x"FF", x"00", x"00", x"EE", x"8A", x"CE", x"8A", x"EA", x"00", x"00", x"FF", x"EE", x"8A", x"CE", x"8A", x"EA", x"FF", x"00", x"00", x"EA", x"8A", x"EE", x"24", x"E4", x"00", x"00", x"FF", x"EA", x"8A", x"EE", x"24", x"E4", x"FF", x"00", x"00", x"FB", x"AA", x"B3", x"AA", x"EA", x"00", x"00", x"FF", x"FB", x"AA", x"B3", x"AA", x"EA", x"FF", x"00", x"00", x"F5", x"95", x"A7", x"C2", x"F2", x"00", x"00", x"FF", x"F5", x"95", x"A7", x"C2", x"F2", x"FF", 
															x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"7F", x"E7", x"C3", x"C3", x"E7", x"7F", x"3F", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"FC", x"FE", x"E7", x"C3", x"C3", x"E7", x"FE", x"FC", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"FC", x"FE", x"E7", x"C3", x"C3", x"E7", x"FE", x"FC", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"01", x"03", x"03", x"07", x"07", x"0F", x"0F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"E0", x"E0", x"F0", x"F0", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"1E", x"3C", x"3C", x"7E", x"7F", x"FF", x"FF", x"FF", x"01", x"03", x"03", x"01", x"00", x"00", x"00", x"00", x"78", x"34", x"34", x"7A", x"FA", x"FD", x"81", x"FF", x"80", x"C8", x"C8", x"84", x"04", x"02", x"7E", x"00", x"0F", x"3F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"FC", x"FC", x"FE", x"FE", x"F8", x"E0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"3F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"60", x"98", x"E6", x"F2", x"0C", x"F0", x"00", x"00", x"80", x"60", x"18", x"0C", x"F0", x"00", x"00", x"00", x"00", x"1C", x"3E", x"36", x"3E", x"1C", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"5A", x"52", x"5A", x"53", x"79", x"00", x"00", x"80", x"DA", x"D2", x"DA", x"D3", x"F9", x"80", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"00", x"00", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"00", x"00", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"00", x"00", x"C0", x"C0", x"00", x"00", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"00", x"00", x"0C", x"0C", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"C0", x"F8", x"C0", x"C0", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"6C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"76", x"14", x"26", x"44", x"76", x"00", x"00", x"01", x"77", x"15", x"27", x"45", x"77", x"01", x"FF", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"C0", x"9C", x"95", x"95", x"D5", x"1D", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"38", x"12", x"52", x"D2", x"D2", x"C2", x"40", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"0A", x"0A", x"AA", x"EA", x"EE", x"E0", x"A0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"E0", x"8E", x"C8", x"8E", x"E2", x"0E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"1E", x"D2", x"D2", x"12", x"D2", x"DE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"04", x"C4", x"C4", x"04", x"C4", x"C4", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"1E", x"C2", x"DE", x"10", x"D0", x"DE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"1E", x"C2", x"CE", x"02", x"C2", x"DE", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"00", x"FF", x"80", x"88", x"88", x"88", x"88", x"88", x"80", x"00", x"00", x"3C", x"04", x"3C", x"20", x"3C", x"00", x"FF", x"80", x"BC", x"84", x"BC", x"A0", x"BC", x"80", x"00", x"00", x"3C", x"04", x"3C", x"04", x"3C", x"00", x"FF", x"80", x"BC", x"84", x"BC", x"84", x"BC", x"80", x"00", x"00", x"0C", x"14", x"24", x"3C", x"04", x"00", x"FF", x"80", x"8C", x"94", x"A4", x"BC", x"84", x"80", x"00", x"00", x"3C", x"20", x"3C", x"04", x"3C", x"00", x"FF", x"80", x"BC", x"A0", x"BC", x"84", x"BC", x"80", 
															x"00", x"00", x"3C", x"20", x"3C", x"24", x"3C", x"00", x"FF", x"80", x"BC", x"A0", x"BC", x"A4", x"BC", x"80", x"00", x"00", x"3C", x"04", x"08", x"10", x"10", x"00", x"FF", x"80", x"BC", x"84", x"88", x"90", x"90", x"80", x"00", x"00", x"3C", x"24", x"3C", x"24", x"3C", x"00", x"FF", x"80", x"BC", x"A4", x"BC", x"A4", x"BC", x"80", x"00", x"00", x"3C", x"24", x"3C", x"04", x"3C", x"00", x"FF", x"80", x"BC", x"A4", x"BC", x"84", x"BC", x"80", x"00", x"00", x"78", x"48", x"48", x"48", x"78", x"00", x"FF", x"01", x"79", x"49", x"49", x"49", x"79", x"01", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"00", x"FF", x"01", x"09", x"09", x"09", x"09", x"09", x"01", x"00", x"00", x"3C", x"04", x"3C", x"20", x"3C", x"00", x"FF", x"01", x"3D", x"05", x"3D", x"21", x"3D", x"01", x"00", x"00", x"3C", x"04", x"3C", x"04", x"3C", x"00", x"FF", x"01", x"3D", x"05", x"3D", x"05", x"3D", x"01", 
															x"00", x"00", x"0C", x"14", x"24", x"3C", x"04", x"00", x"FF", x"01", x"0D", x"15", x"25", x"3D", x"05", x"01", x"00", x"00", x"3C", x"20", x"3C", x"04", x"3C", x"00", x"FF", x"01", x"3D", x"21", x"3D", x"05", x"3D", x"01", x"00", x"00", x"3C", x"20", x"3C", x"24", x"3C", x"00", x"FF", x"01", x"3D", x"21", x"3D", x"25", x"3D", x"01", x"00", x"00", x"3C", x"04", x"08", x"10", x"10", x"00", x"FF", x"01", x"3D", x"05", x"09", x"11", x"11", x"01", x"00", x"00", x"3C", x"24", x"3C", x"24", x"3C", x"00", x"FF", x"01", x"3D", x"25", x"3D", x"25", x"3D", x"01", x"00", x"00", x"3C", x"24", x"3C", x"04", x"3C", x"00", x"FF", x"01", x"3D", x"25", x"3D", x"05", x"3D", x"01", x"00", x"B4", x"A4", x"B4", x"A4", x"36", x"00", x"00", x"01", x"B5", x"A5", x"B5", x"A5", x"37", x"01", x"FF", x"00", x"57", x"75", x"77", x"55", x"55", x"00", x"00", x"80", x"D7", x"F5", x"F7", x"D5", x"D5", x"80", x"FF");
	
	constant GAME_1942_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"58", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"06", x"1C", x"30", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"06", x"1C", x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"60", x"7C", x"66", x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"60", x"7C", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"06", x"0C", x"18", x"30", x"30", x"30", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"3C", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"3E", x"06", x"04", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C0", x"C0", x"C0", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C0", x"C0", x"CE", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"CC", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"CC", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"D6", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"DE", x"CE", x"C6", x"C6", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"CE", x"C6", x"FC", x"D8", x"CC", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"66", x"66", x"24", x"18", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"D6", x"FE", x"6C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"44", x"6C", x"38", x"38", x"6C", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"06", x"0C", x"18", x"30", x"60", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"CE", x"DC", x"38", x"76", x"E6", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"40", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"D8", x"CC", x"C6", x"00", x"FE", x"FF", x"E7", x"FF", x"FE", x"EF", x"E7", x"63", 
															x"01", x"03", x"0F", x"1B", x"37", x"27", x"73", x"79", x"00", x"02", x"0C", x"1C", x"38", x"38", x"7C", x"7E", x"00", x"C0", x"70", x"38", x"1C", x"3C", x"7E", x"FF", x"00", x"C0", x"F0", x"F8", x"FC", x"CC", x"82", x"00", x"FF", x"7F", x"3E", x"3E", x"1D", x"0F", x"03", x"00", x"00", x"41", x"33", x"3F", x"1F", x"0F", x"03", x"00", x"FE", x"EE", x"F4", x"FC", x"F8", x"F0", x"C0", x"80", x"7E", x"3E", x"1C", x"1C", x"38", x"30", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"22", x"02", x"3E", x"22", x"2A", x"2A", x"23", x"FE", x"EE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"08", x"08", x"08", x"58", x"F0", x"00", x"00", x"00", x"58", x"58", x"F8", x"F8", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"32", 
															x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"18", x"18", x"00", x"00", x"18", x"18", x"18", x"18", x"00", x"00", x"18", x"18", x"18", x"18", x"18", x"18", x"06", x"C6", x"C0", x"00", x"06", x"C6", x"C6", x"C0", x"00", x"00", x"06", x"C6", x"C6", x"C6", x"C6", x"C0", x"00", x"02", x"05", x"05", x"00", x"00", x"65", x"1D", x"00", x"1F", x"07", x"07", x"7F", x"FF", x"7F", x"1F", x"10", x"38", x"19", x"19", x"11", x"00", x"C7", x"EF", x"10", x"FF", x"29", x"29", x"EF", x"FF", x"FF", x"FF", x"7F", x"20", x"00", x"10", x"00", x"10", x"5F", x"00", x"5F", x"00", x"70", x"70", x"20", x"7F", x"FF", x"20", x"FC", x"08", x"00", x"04", x"00", x"04", x"F6", x"00", x"F4", x"00", x"1C", x"1C", x"08", x"FC", x"FE", x"08", x"02", x"02", x"05", x"05", x"7F", x"1F", x"03", x"01", x"00", x"05", x"07", x"FF", x"7F", x"1F", x"03", x"01", 
															x"00", x"08", x"19", x"39", x"FF", x"FF", x"01", x"83", x"10", x"39", x"29", x"EF", x"EF", x"FF", x"01", x"83", x"82", x"FF", x"C6", x"44", x"00", x"00", x"00", x"00", x"82", x"FF", x"C6", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"02", x"00", x"00", x"00", x"02", x"07", x"7F", x"07", x"02", x"00", x"00", x"00", x"00", x"01", x"29", x"6D", x"D6", x"44", x"00", x"00", x"38", x"7D", x"FF", x"55", x"D6", x"44", x"00", x"00", x"00", x"00", x"00", x"08", x"22", x"42", x"40", x"00", x"00", x"00", x"44", x"6C", x"FF", x"C6", x"C6", x"00", x"0C", x"04", x"09", x"03", x"0E", x"0C", x"00", x"03", x"0F", x"7F", x"FF", x"07", x"0A", x"08", x"00", x"00", x"92", x"8A", x"2D", x"09", x"28", x"38", x"10", x"FF", x"FF", x"FF", x"FF", x"39", x"38", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"50", x"58", x"5F", x"00", x"00", x"00", x"00", x"20", x"FF", x"FF", x"FF", 
															x"02", x"0C", x"01", x"01", x"01", x"00", x"02", x"01", x"03", x"0F", x"3E", x"7E", x"3E", x"03", x"03", x"0F", x"40", x"30", x"AC", x"A0", x"A0", x"00", x"40", x"80", x"C0", x"F0", x"7C", x"7E", x"7C", x"C0", x"C0", x"F0", x"00", x"00", x"00", x"0C", x"08", x"08", x"00", x"00", x"00", x"00", x"10", x"FE", x"7C", x"38", x"10", x"10", x"00", x"02", x"0F", x"21", x"00", x"01", x"02", x"01", x"01", x"03", x"0E", x"3E", x"7F", x"03", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"2C", x"00", x"00", x"00", x"00", x"00", x"10", x"FE", x"7C", x"00", x"00", x"00", x"02", x"01", x"01", x"02", x"03", x"00", x"01", x"01", x"0F", x"00", x"02", x"7F", x"03", x"01", x"02", x"01", x"00", x"04", x"00", x"00", x"00", x"01", x"03", x"03", x"7F", x"3F", x"0F", x"03", x"01", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"FE", x"10", x"00", x"00", x"00", x"00", x"00", 
															x"01", x"02", x"00", x"00", x"04", x"00", x"00", x"00", x"0F", x"03", x"03", x"3F", x"7F", x"3F", x"0F", x"07", x"28", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"38", x"10", x"38", x"7C", x"FE", x"10", x"00", x"00", x"04", x"08", x"16", x"32", x"16", x"00", x"02", x"01", x"07", x"0F", x"1D", x"3D", x"1D", x"03", x"03", x"0F", x"80", x"A0", x"00", x"80", x"80", x"80", x"80", x"00", x"C0", x"E0", x"F8", x"FC", x"F8", x"80", x"80", x"E0", x"00", x"10", x"80", x"00", x"B8", x"10", x"00", x"00", x"08", x"18", x"B8", x"FC", x"B8", x"18", x"08", x"00", x"28", x"60", x"48", x"40", x"28", x"28", x"10", x"00", x"38", x"38", x"38", x"38", x"38", x"38", x"FE", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"00", x"08", x"00", x"00", x"10", x"F0", x"70", x"30", x"10", x"18", x"00", x"00", x"00", x"02", x"00", x"00", x"02", x"01", x"03", x"0F", x"3F", x"7F", x"3F", x"03", x"03", x"0F", 
															x"C0", x"20", x"10", x"58", x"30", x"80", x"80", x"40", x"C0", x"E0", x"F0", x"F8", x"F8", x"80", x"80", x"E0", x"00", x"00", x"00", x"0C", x"08", x"08", x"00", x"28", x"00", x"00", x"10", x"FC", x"7C", x"38", x"10", x"38", x"00", x"08", x"10", x"10", x"20", x"20", x"42", x"35", x"00", x"08", x"18", x"18", x"38", x"38", x"7E", x"CF", x"00", x"00", x"02", x"03", x"00", x"03", x"02", x"00", x"00", x"02", x"03", x"03", x"07", x"03", x"03", x"02", x"00", x"02", x"02", x"02", x"02", x"02", x"13", x"0D", x"00", x"02", x"02", x"02", x"12", x"12", x"17", x"73", x"00", x"00", x"00", x"00", x"00", x"08", x"40", x"A0", x"00", x"10", x"18", x"18", x"1C", x"1C", x"7C", x"FE", x"00", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"40", x"C0", x"C0", x"E0", x"C0", x"C0", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"40", x"80", x"00", x"08", x"1C", x"1C", x"9E", x"9F", x"FF", x"FF", 
															x"00", x"00", x"00", x"80", x"00", x"B8", x"10", x"00", x"00", x"08", x"18", x"B8", x"FC", x"B8", x"18", x"08", x"00", x"00", x"00", x"04", x"04", x"02", x"02", x"41", x"00", x"00", x"08", x"1C", x"1C", x"9E", x"9E", x"FF", x"9C", x"71", x"1E", x"02", x"04", x"04", x"00", x"00", x"E3", x"FF", x"9E", x"9E", x"1C", x"1C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"10", x"00", x"00", x"10", x"30", x"70", x"F8", x"70", x"30", x"10", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"03", x"03", x"03", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"18", x"58", x"A0", x"50", x"20", x"00", x"20", x"90", x"D8", x"EC", x"D2", x"B8", x"FC", x"00", x"18", x"08", x"06", x"02", x"00", x"00", x"00", x"1D", x"1E", x"0F", x"0F", x"03", x"00", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"08", x"1C", x"02", x"15", x"5C", x"80", x"00", x"00", x"08", x"1C", x"9E", x"9F", x"E3", x"FF", x"7B", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"FF", x"9F", x"9E", x"1C", x"1C", x"08", x"00", x"00", x"02", x"00", x"02", x"00", x"14", x"04", x"00", x"02", x"03", x"01", x"03", x"03", x"1E", x"1E", x"0F", x"03", x"00", x"0E", x"33", x"40", x"35", x"00", x"00", x"00", x"40", x"40", x"7F", x"7F", x"7F", x"40", x"40", x"00", x"00", x"00", x"30", x"00", x"80", x"00", x"00", x"00", x"08", x"18", x"38", x"FC", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"48", x"80", x"00", x"08", x"1C", x"1C", x"9E", x"9E", x"FF", x"FF", x"61", x"89", x"12", x"1C", x"08", x"00", x"00", x"00", x"FF", x"9F", x"9E", x"1C", x"18", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"B8", x"08", x"00", x"00", x"08", x"18", x"B8", x"FC", x"B8", x"18", x"00", x"00", 
															x"00", x"00", x"01", x"01", x"0C", x"08", x"01", x"33", x"00", x"06", x"0F", x"1F", x"33", x"77", x"7F", x"3E", x"00", x"00", x"80", x"80", x"34", x"3A", x"B6", x"DC", x"00", x"60", x"F0", x"F8", x"CC", x"EE", x"FE", x"7C", x"33", x"03", x"2D", x"1E", x"17", x"0F", x"06", x"00", x"3E", x"7F", x"77", x"33", x"1F", x"0F", x"06", x"00", x"EC", x"DE", x"FE", x"FC", x"F8", x"F0", x"60", x"00", x"7C", x"FE", x"EE", x"CC", x"F8", x"F0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"CC", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"CC", x"FC", x"C0", x"DD", x"D5", x"D5", x"DC", x"00", x"EE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"10", x"50", x"50", x"F0", x"A0", x"00", x"00", x"00", x"10", x"58", x"58", x"F8", x"F8", x"F0", x"EE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"22", x"02", x"3E", x"22", x"2A", x"2A", x"23", x"FE", 
															x"00", x"00", x"10", x"00", x"08", x"10", x"1C", x"14", x"00", x"00", x"10", x"10", x"38", x"28", x"6C", x"EE", x"00", x"00", x"54", x"00", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"03", x"03", x"01", x"01", x"00", x"C0", x"40", x"D4", x"00", x"80", x"00", x"00", x"00", x"F8", x"FC", x"FC", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"20", x"03", x"06", x"00", x"00", x"00", x"00", x"78", x"7E", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"20", x"40", x"80", x"00", x"00", x"00", x"00", x"30", x"50", x"A0", x"40", x"04", x"00", x"09", x"04", x"00", x"00", x"00", x"00", x"07", x"07", x"0F", x"1C", x"18", x"00", x"00", x"00", x"40", x"C0", x"80", x"00", x"10", x"20", x"00", x"00", x"C0", x"E0", x"E0", x"F0", x"70", x"30", x"30", x"00", x"00", x"00", x"00", x"E4", x"50", x"C0", x"00", x"00", x"80", x"C0", x"F0", x"1C", x"F0", x"C0", x"80", x"00", 
															x"00", x"04", x"00", x"04", x"00", x"04", x"00", x"00", x"00", x"06", x"07", x"07", x"07", x"07", x"1F", x"7F", x"15", x"07", x"00", x"04", x"00", x"04", x"00", x"00", x"1F", x"07", x"07", x"07", x"07", x"06", x"00", x"00", x"24", x"08", x"28", x"08", x"28", x"10", x"00", x"00", x"FE", x"70", x"70", x"30", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"02", x"00", x"00", x"01", x"01", x"01", x"03", x"3F", x"3F", x"1F", x"00", x"00", x"40", x"80", x"00", x"A0", x"50", x"60", x"00", x"C0", x"C0", x"80", x"00", x"F0", x"F0", x"F0", x"04", x"0C", x"44", x"08", x"20", x"10", x"00", x"00", x"78", x"78", x"78", x"38", x"38", x"10", x"00", x"00", x"00", x"00", x"04", x"08", x"20", x"10", x"40", x"08", x"00", x"1C", x"1C", x"18", x"30", x"30", x"70", x"78", x"48", x"14", x"0C", x"14", x"08", x"10", x"00", x"00", x"7E", x"38", x"38", x"38", x"38", x"10", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"16", x"0C", x"05", x"00", x"01", x"01", x"01", x"01", x"1F", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"C0", x"C0", x"80", x"00", x"FC", x"FC", x"F8", x"0C", x"04", x"08", x"00", x"08", x"00", x"00", x"00", x"FE", x"7C", x"38", x"38", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"07", x"7F", x"7F", x"3F", x"00", x"00", x"80", x"00", x"C0", x"40", x"C0", x"40", x"00", x"00", x"80", x"80", x"C0", x"FC", x"FC", x"F8", x"00", x"01", x"00", x"10", x"00", x"01", x"05", x"01", x"00", x"01", x"01", x"33", x"33", x"3E", x"FE", x"FE", x"00", x"00", x"00", x"88", x"00", x"E0", x"40", x"C0", x"00", x"00", x"00", x"98", x"98", x"F8", x"FE", x"FE", x"04", x"02", x"00", x"20", x"02", x"00", x"00", x"00", x"7F", x"33", x"31", x"01", x"0F", x"1F", x"0D", x"00", 
															x"60", x"80", x"00", x"08", x"C0", x"80", x"00", x"00", x"FC", x"98", x"18", x"00", x"E0", x"F0", x"60", x"00", x"00", x"00", x"01", x"22", x"00", x"05", x"2B", x"02", x"00", x"03", x"37", x"3E", x"1F", x"3F", x"1B", x"03", x"00", x"00", x"00", x"00", x"00", x"A0", x"40", x"A0", x"00", x"00", x"00", x"18", x"78", x"D0", x"B0", x"60", x"00", x"04", x"12", x"20", x"24", x"18", x"00", x"00", x"03", x"E7", x"FE", x"7C", x"3C", x"1E", x"0E", x"06", x"64", x"C8", x"20", x"40", x"00", x"48", x"00", x"00", x"F6", x"FE", x"3C", x"78", x"7C", x"2C", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"11", x"02", x"00", x"00", x"01", x"07", x"27", x"71", x"71", x"33", x"7F", x"00", x"00", x"00", x"08", x"00", x"40", x"00", x"E2", x"C0", x"C0", x"F8", x"F8", x"E0", x"E0", x"F8", x"1E", x"32", x"11", x"01", x"00", x"08", x"00", x"00", x"00", x"33", x"71", x"71", x"27", x"07", x"01", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"20", x"51", x"01", x"4D", x"00", x"00", x"01", x"03", x"FB", x"72", x"72", x"FE", x"00", x"00", x"00", x"00", x"88", x"14", x"80", x"52", x"00", x"00", x"00", x"80", x"BE", x"9C", x"9C", x"FF", x"08", x"54", x"18", x"55", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"7E", x"26", x"03", x"03", x"03", x"E2", x"54", x"E4", x"74", x"C0", x"00", x"80", x"00", x"FF", x"FF", x"FF", x"FC", x"C8", x"80", x"80", x"80", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"01", x"03", x"0F", x"3F", x"1F", x"01", x"00", x"80", x"00", x"80", x"C0", x"80", x"80", x"00", x"00", x"80", x"00", x"80", x"E0", x"F8", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"0F", x"01", x"00", x"00", x"A0", x"10", x"20", x"80", x"00", x"28", x"E4", x"90", x"F0", x"F0", x"F0", x"94", x"84", x"FC", x"1C", 
															x"A8", x"80", x"00", x"A0", x"10", x"20", x"80", x"00", x"FC", x"84", x"94", x"F0", x"F0", x"F0", x"90", x"80", x"00", x"02", x"00", x"0D", x"03", x"08", x"00", x"18", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"FF", x"E7", x"AA", x"0F", x"0C", x"0A", x"00", x"06", x"03", x"00", x"FF", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"38", x"38", x"3C", x"3D", x"7F", x"3D", x"30", x"20", x"00", x"00", x"00", x"00", x"00", x"3D", x"3C", x"38", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"38", x"38", x"78", x"E0", x"90", x"48", x"45", x"26", x"28", x"11", x"02", x"E0", x"F1", x"78", x"7D", x"3F", x"3F", x"1F", x"1F", x"28", x"90", x"18", x"24", x"42", x"31", x"0D", x"03", x"FA", x"F0", x"F8", x"FC", x"FE", x"3F", x"0F", x"03", 
															x"00", x"80", x"8C", x"34", x"48", x"28", x"50", x"A6", x"80", x"C0", x"AC", x"3C", x"78", x"DC", x"B2", x"67", x"31", x"12", x"20", x"18", x"3B", x"55", x"A0", x"40", x"3E", x"1D", x"3F", x"37", x"2F", x"7D", x"E0", x"C0", x"62", x"55", x"4A", x"14", x"0A", x"01", x"07", x"00", x"63", x"77", x"7E", x"3C", x"1E", x"2F", x"07", x"00", x"1E", x"16", x"06", x"0C", x"06", x"16", x"16", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"0E", x"16", x"16", x"16", x"1E", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"10", x"10", x"1E", x"06", x"06", x"16", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"16", x"10", x"1E", x"16", x"16", x"16", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"16", x"06", x"06", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"1E", x"16", x"16", x"1C", x"16", x"16", x"16", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"16", x"16", x"16", x"1E", x"06", x"0C", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"16", x"06", x"08", x"10", x"16", x"16", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"AA", x"AA", x"AA", x"AA", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"80", x"8E", x"EA", x"2A", x"2A", x"AA", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"A0", x"A0", x"A0", x"A0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A8", x"E0", x"20", x"00", x"08", x"00", x"00", x"00", x"F8", x"E0", x"E0", x"F8", x"F8", x"C0", x"C0", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"6C", x"04", x"28", x"04", x"14", x"00", x"10", x"FF", x"7C", x"7C", x"38", x"7C", x"6C", x"00", x"00", x"00", x"05", x"00", x"00", x"00", x"00", x"7F", x"FF", x"7F", x"0F", x"00", x"00", x"00", x"00", x"3E", x"3C", x"06", x"07", x"C6", x"7C", x"54", x"00", x"C7", x"C7", x"FF", x"FF", x"FE", x"44", x"6C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"05", x"38", x"38", x"38", x"10", x"38", x"FE", x"FF", x"D7", x"00", x"00", x"01", x"02", x"12", x"21", x"01", x"02", x"00", x"00", x"0F", x"03", x"FF", x"32", x"32", x"35", x"00", x"00", x"00", x"80", x"90", x"08", x"00", x"C0", x"00", x"00", x"E0", x"80", x"FE", x"98", x"98", x"58", 
															x"00", x"00", x"00", x"05", x"01", x"00", x"00", x"00", x"7F", x"FF", x"7F", x"0F", x"01", x"00", x"00", x"00", x"2C", x"04", x"06", x"17", x"97", x"44", x"00", x"00", x"D7", x"FF", x"FF", x"EF", x"EF", x"7C", x"38", x"38", x"00", x"00", x"00", x"10", x"00", x"00", x"00", x"00", x"03", x"01", x"23", x"3F", x"2F", x"23", x"01", x"00", x"80", x"00", x"80", x"50", x"00", x"80", x"00", x"00", x"80", x"00", x"88", x"F8", x"E8", x"88", x"00", x"00", x"00", x"40", x"A0", x"20", x"11", x"20", x"41", x"04", x"00", x"F0", x"E0", x"E0", x"FF", x"FF", x"FF", x"FC", x"00", x"00", x"02", x"05", x"08", x"04", x"0B", x"00", x"00", x"00", x"0F", x"07", x"7F", x"FF", x"3F", x"01", x"00", x"00", x"10", x"10", x"84", x"46", x"55", x"24", x"10", x"38", x"AB", x"29", x"FF", x"FF", x"FF", x"FF", x"24", x"10", x"20", x"00", x"00", x"28", x"84", x"10", x"FE", x"28", x"38", x"10", x"10", x"7C", x"D6", x"00", 
															x"10", x"54", x"54", x"04", x"54", x"04", x"04", x"3C", x"28", x"28", x"28", x"7C", x"28", x"7C", x"7C", x"44", x"7C", x"4C", x"04", x"0C", x"04", x"0E", x"06", x"0E", x"00", x"38", x"7C", x"7C", x"7F", x"7F", x"7F", x"7F", x"07", x"87", x"07", x"AF", x"3F", x"97", x"06", x"04", x"FF", x"FF", x"FF", x"D7", x"C7", x"EF", x"FE", x"7C", x"82", x"82", x"86", x"04", x"00", x"00", x"00", x"00", x"7C", x"7C", x"7C", x"7C", x"38", x"38", x"38", x"38", x"00", x"00", x"00", x"00", x"0A", x"03", x"03", x"01", x"07", x"3F", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"80", x"80", x"00", x"C0", x"F8", x"FE", x"FF", x"FE", x"00", x"00", x"00", x"00", x"10", x"28", x"00", x"00", x"08", x"08", x"10", x"10", x"FE", x"38", x"38", x"38", x"38", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"07", x"01", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"0A", x"01", x"00", x"7F", x"FF", x"FF", x"FF", x"FF", x"1F", x"01", x"00", x"00", x"00", x"00", x"AA", x"55", x"0A", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"1F", x"03", x"01", x"00", x"00", x"80", x"95", x"EA", x"D0", x"C0", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"C0", x"80", x"10", x"10", x"00", x"10", x"38", x"28", x"00", x"00", x"00", x"28", x"38", x"28", x"00", x"11", x"38", x"38", x"10", x"20", x"43", x"84", x"28", x"18", x"20", x"00", x"FF", x"FF", x"FF", x"FF", x"10", x"38", x"38", x"38", x"44", x"4C", x"00", x"00", x"08", x"2C", x"BA", x"10", x"38", x"38", x"10", x"10", x"7C", x"FE", x"82", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"01", x"00", x"00", x"04", x"0A", x"02", x"01", x"02", x"34", x"40", x"00", x"1F", x"0E", x"0E", x"FF", x"FF", x"FF", x"7F", 
															x"40", x"28", x"5C", x"8C", x"16", x"22", x"23", x"F5", x"40", x"28", x"5C", x"8C", x"1E", x"3F", x"3F", x"FB", x"17", x"3B", x"4B", x"A4", x"3A", x"53", x"91", x"21", x"18", x"3C", x"4C", x"A7", x"3B", x"53", x"91", x"21", x"82", x"49", x"E4", x"7C", x"2D", x"21", x"4F", x"07", x"82", x"49", x"E5", x"7F", x"3E", x"3E", x"70", x"38", x"CF", x"4D", x"23", x"73", x"3B", x"30", x"60", x"C0", x"F0", x"72", x"3C", x"7C", x"3C", x"3F", x"66", x"C0", x"22", x"04", x"08", x"64", x"C2", x"83", x"07", x"05", x"00", x"00", x"08", x"04", x"02", x"03", x"07", x"07", x"38", x"24", x"04", x"4F", x"DB", x"B1", x"2D", x"EF", x"00", x"04", x"04", x"4F", x"DF", x"FF", x"F3", x"F1", x"12", x"8A", x"14", x"79", x"17", x"D3", x"41", x"0A", x"15", x"0D", x"1B", x"7F", x"1F", x"1F", x"0F", x"0D", x"D5", x"9B", x"AF", x"66", x"9C", x"FA", x"F5", x"65", x"FB", x"FF", x"DF", x"9F", x"FF", x"FD", x"FB", x"FB", 
															x"15", x"06", x"43", x"65", x"28", x"06", x"01", x"00", x"16", x"07", x"03", x"05", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"09", x"04", x"03", x"02", x"10", x"00", x"00", x"22", x"49", x"44", x"03", x"00", x"00", x"00", x"14", x"58", x"2C", x"E6", x"C7", x"20", x"82", x"10", x"14", x"58", x"3C", x"FE", x"FF", x"06", x"0C", x"08", x"5D", x"3F", x"0C", x"04", x"0A", x"07", x"8F", x"0F", x"5F", x"3F", x"8F", x"47", x"8B", x"84", x"CC", x"D2", x"E1", x"F9", x"6E", x"62", x"42", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"0E", x"0D", x"10", x"00", x"00", x"00", x"00", x"07", x"2E", x"0D", x"90", x"02", x"40", x"20", x"04", x"00", x"00", x"00", x"00", x"00", x"02", x"01", x"02", x"22", x"40", x"09", x"40", x"20", x"02", x"81", x"23", x"00", x"00", x"00", x"08", x"10", x"20", x"C0", x"60", x"09", x"40", x"02", x"48", x"10", x"24", x"C0", x"E2", 
															x"00", x"00", x"01", x"17", x"0F", x"0F", x"1E", x"3C", x"00", x"00", x"01", x"17", x"0F", x"0F", x"1F", x"3F", x"00", x"00", x"C2", x"EC", x"F8", x"70", x"58", x"3C", x"00", x"00", x"C2", x"EC", x"F8", x"F0", x"F8", x"FC", x"00", x"09", x"07", x"5F", x"3C", x"38", x"70", x"60", x"00", x"09", x"07", x"5F", x"3F", x"3F", x"7F", x"7F", x"40", x"E0", x"FA", x"BC", x"3E", x"1E", x"1F", x"0F", x"40", x"E0", x"FA", x"FC", x"FE", x"FE", x"FF", x"FF", x"00", x"13", x"0E", x"B8", x"61", x"61", x"C3", x"C7", x"00", x"13", x"0F", x"BF", x"7E", x"7E", x"FC", x"F8", x"80", x"E4", x"38", x"1C", x"06", x"82", x"C3", x"E3", x"80", x"E4", x"F8", x"FC", x"FE", x"7E", x"3F", x"1F", x"01", x"04", x"10", x"48", x"21", x"03", x"87", x"03", x"01", x"04", x"11", x"4A", x"24", x"48", x"80", x"28", x"00", x"50", x"08", x"21", x"42", x"E0", x"E0", x"F5", x"00", x"50", x"48", x"A1", x"12", x"04", x"0A", x"05", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"7F", x"7F", x"FF", x"FF", x"00", x"00", x"03", x"0E", x"18", x"10", x"30", x"20", x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"00", x"03", x"0F", x"0E", x"1C", x"18", x"00", x"00", x"00", x"03", x"0F", x"0F", x"1F", x"1F", x"00", x"00", x"00", x"00", x"03", x"07", x"0E", x"0C", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"0F", x"00", x"3C", x"7E", x"FF", x"FF", x"7E", x"3C", x"00", x"00", x"3C", x"7E", x"FF", x"FF", x"7E", x"3C", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"18", x"00", x"00", x"00", x"A0", x"C0", x"E0", x"C0", x"E0", x"C0", x"E0", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"58", x"58", x"F8", x"F8", x"F0", x"00", x"00", x"00", x"08", x"08", x"08", x"58", x"F0", 
															x"00", x"00", x"00", x"00", x"00", x"14", x"16", x"F6", x"00", x"00", x"00", x"00", x"08", x"FE", x"FF", x"FE", x"00", x"00", x"10", x"08", x"08", x"10", x"16", x"18", x"20", x"20", x"70", x"F8", x"F8", x"70", x"77", x"FF", x"00", x"00", x"04", x"02", x"02", x"04", x"04", x"06", x"08", x"08", x"1C", x"3E", x"3E", x"1C", x"DC", x"FF", x"E1", x"01", x"03", x"01", x"05", x"02", x"00", x"00", x"FF", x"FF", x"FF", x"07", x"07", x"0F", x"00", x"00", x"8C", x"8C", x"8E", x"08", x"08", x"08", x"28", x"10", x"FF", x"FF", x"FF", x"39", x"39", x"BB", x"38", x"10", x"6E", x"60", x"70", x"40", x"40", x"80", x"00", x"00", x"FE", x"FF", x"FE", x"C0", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"28", x"2C", x"00", x"28", x"00", x"00", x"10", x"10", x"7F", x"3F", x"10", x"38", x"10", x"02", x"22", x"FE", x"FF", x"03", x"01", x"00", x"00", x"0F", x"3F", x"FF", x"FF", x"03", x"01", x"00", x"00", 
															x"C8", x"88", x"CC", x"FF", x"BB", x"39", x"38", x"10", x"FF", x"FF", x"FF", x"FF", x"BB", x"39", x"38", x"10", x"00", x"00", x"02", x"00", x"7F", x"01", x"00", x"00", x"01", x"01", x"07", x"01", x"7F", x"01", x"00", x"00", x"00", x"10", x"9A", x"8A", x"EF", x"BB", x"38", x"00", x"01", x"01", x"FF", x"BB", x"EF", x"BB", x"38", x"00", x"00", x"00", x"04", x"24", x"04", x"04", x"01", x"01", x"01", x"03", x"7F", x"3F", x"0F", x"07", x"03", x"03", x"82", x"00", x"92", x"10", x"82", x"00", x"83", x"01", x"93", x"BB", x"EF", x"EF", x"FF", x"83", x"83", x"01", x"48", x"90", x"10", x"00", x"00", x"00", x"00", x"00", x"7F", x"FF", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"80", x"74", x"0F", x"00", x"17", x"08", x"01", x"0A", x"FF", x"7F", x"07", x"08", x"1F", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"58", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"06", x"1C", x"30", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"06", x"1C", x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"1E", x"36", x"66", x"7F", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"60", x"7C", x"66", x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"60", x"7C", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"06", x"0C", x"18", x"30", x"30", x"30", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"3C", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"3E", x"06", x"04", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C0", x"C0", x"C0", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FE", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"D6", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"CE", x"C6", x"FC", x"D8", x"CC", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"44", x"9A", x"A2", x"9A", x"44", x"38", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"18", x"18", x"18", x"18", x"18", x"18", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CF", x"87", x"13", x"4B", x"BF", x"FF", x"FF", x"FF", x"30", x"78", x"FC", x"FC", x"70", x"18", x"3C", x"18", x"01", x"F9", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"07", x"07", x"07", x"1F", x"1F", x"1F", x"11", x"01", x"02", x"1A", x"1A", x"02", x"3E", x"3E", x"1F", x"0F", x"3E", x"26", x"26", x"3E", x"3E", x"3E", x"14", x"79", x"CB", x"35", x"51", x"0A", x"D6", x"31", x"FF", x"CF", x"BF", x"FF", x"FF", x"FF", x"FF", x"FF", x"02", x"CF", x"FF", x"FB", x"B9", x"EF", x"FF", x"FF", x"FD", x"38", x"42", x"04", x"47", x"12", x"08", x"00", x"0D", x"CD", x"CC", x"D9", x"F3", x"E6", x"FC", x"F8", x"FF", x"7F", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", 
															x"23", x"57", x"6A", x"11", x"2A", x"76", x"83", x"70", x"DC", x"E9", x"F7", x"EF", x"DD", x"BF", x"FF", x"FF", x"45", x"2B", x"56", x"0C", x"14", x"FD", x"C1", x"06", x"BB", x"D7", x"EF", x"F7", x"FB", x"77", x"FF", x"FF", x"00", x"00", x"00", x"01", x"07", x"1C", x"70", x"C0", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", x"07", x"1C", x"70", x"CF", x"0F", x"6F", x"6F", x"6F", x"00", x"03", x"0F", x"3F", x"F8", x"98", x"9F", x"FF", x"E0", x"38", x"0E", x"F3", x"F0", x"F6", x"F6", x"F6", x"00", x"C0", x"F0", x"FC", x"1F", x"19", x"F9", x"FF", x"00", x"00", x"00", x"80", x"E0", x"38", x"0E", x"03", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"80", x"00", x"80", x"00", x"80", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", 
															x"00", x"04", x"00", x"04", x"00", x"04", x"00", x"04", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"20", x"00", x"20", x"00", x"20", x"00", x"20", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"10", x"00", x"10", x"00", x"10", x"00", x"10", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"08", x"00", x"08", x"00", x"08", x"00", x"08", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"40", x"00", x"40", x"00", x"40", x"00", x"40", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"02", x"00", x"02", x"00", x"02", x"00", x"02", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"DE", x"CE", x"C6", x"C6", 
															x"FF", x"FF", x"FF", x"1C", x"1C", x"1C", x"1C", x"1C", x"00", x"00", x"00", x"E3", x"E3", x"E3", x"E3", x"E3", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"E3", x"E3", x"E3", x"E3", x"E3", x"E3", x"E3", x"E3", x"00", x"00", x"0F", x"1F", x"3C", x"38", x"30", x"30", x"FF", x"F0", x"E0", x"C0", x"80", x"83", x"87", x"87", x"00", x"00", x"F0", x"F8", x"3C", x"1C", x"0C", x"0C", x"FF", x"0F", x"07", x"03", x"01", x"C1", x"E1", x"E1", x"38", x"1C", x"0F", x"07", x"0F", x"1C", x"38", x"30", x"83", x"C0", x"E0", x"F0", x"E0", x"C0", x"83", x"87", x"1C", x"38", x"F0", x"E0", x"F0", x"38", x"1C", x"0C", x"C1", x"03", x"07", x"0F", x"07", x"03", x"C1", x"E1", x"30", x"30", x"38", x"3C", x"1F", x"0F", x"00", x"00", x"87", x"87", x"83", x"80", x"C0", x"E0", x"F0", x"FF", 
															x"0C", x"0C", x"1C", x"3C", x"F8", x"F0", x"00", x"00", x"E1", x"E1", x"C1", x"01", x"03", x"07", x"0F", x"FF", x"1F", x"70", x"C1", x"FB", x"F8", x"FA", x"F9", x"C8", x"E0", x"8F", x"3E", x"04", x"07", x"07", x"7F", x"7F", x"EF", x"EC", x"EE", x"4E", x"78", x"49", x"7A", x"FF", x"10", x"5B", x"59", x"F9", x"FF", x"FF", x"FF", x"FF", x"FC", x"06", x"13", x"89", x"85", x"C7", x"67", x"37", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A0", x"81", x"F9", x"F9", x"F9", x"F9", x"CB", x"A2", x"7F", x"7E", x"06", x"06", x"06", x"7E", x"7E", x"7F", x"F8", x"FC", x"F9", x"F1", x"E9", x"C5", x"46", x"BD", x"07", x"47", x"2F", x"1F", x"3F", x"FF", x"FF", x"FF", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"83", x"8F", x"3F", x"E6", x"E4", x"F8", x"F0", x"41", x"7F", x"7E", x"C4", x"DD", x"9F", x"3F", x"8F", x"BF", 
															x"FF", x"00", x"FC", x"02", x"39", x"7C", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C7", x"93", x"39", x"26", x"CC", x"38", x"18", x"0C", x"86", x"43", x"23", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C1", x"73", x"F3", x"53", x"C3", x"43", x"F3", x"73", x"BF", x"8E", x"BE", x"BE", x"BE", x"BE", x"8E", x"BE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7D", x"7C", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"23", x"A3", x"A3", x"A3", x"A3", x"BF", x"BF", x"BF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"FF", x"F1", x"73", x"D3", x"43", x"F3", x"73", x"D3", x"43", x"8F", x"BE", x"BE", x"BE", x"8E", x"BE", x"BE", x"BE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"7C", x"7D", x"A3", x"A3", x"BF", x"BF", x"BF", x"A3", x"A3", x"BF", x"FF", x"FF", x"E7", x"E7", x"FF", x"FF", x"FF", x"E7", 
															x"E1", x"BC", x"A6", x"E6", x"BC", x"A6", x"E7", x"9D", x"BF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"7F", x"3E", x"1C", x"00", x"29", x"83", x"39", x"93", x"C7", x"FF", x"FF", x"FF", x"D7", x"FF", x"A7", x"BF", x"2F", x"6F", x"CF", x"9F", x"FF", x"3D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"84", x"B4", x"B5", x"85", x"84", x"BC", x"A2", x"A3", x"7B", x"CB", x"4A", x"7B", x"7B", x"47", x"5F", x"5F", x"FE", x"00", x"80", x"FC", x"7C", x"7C", x"01", x"FF", x"FF", x"FF", x"FF", x"87", x"87", x"FF", x"FF", x"FF", x"1D", x"1D", x"1D", x"3D", x"6C", x"CD", x"8D", x"0D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AB", x"A3", x"97", x"C4", x"40", x"77", x"37", x"1F", x"56", x"56", x"E7", x"F7", x"F7", x"F7", x"F7", x"FF", x"C0", x"C1", x"C1", x"0F", x"0F", x"FF", x"FF", x"FF", x"7F", x"7E", x"FF", x"F2", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"02", x"20", x"00", x"04", x"40", x"92", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"2C", x"FE", x"00", x"08", x"40", x"10", x"02", x"40", x"82", x"00", x"00", x"00", x"00", x"00", x"08", x"1C", x"7C", x"FF", x"10", x"00", x"04", x"40", x"01", x"92", x"30", x"40", x"00", x"00", x"00", x"00", x"00", x"09", x"1F", x"3F", x"10", x"A4", x"00", x"52", x"20", x"00", x"08", x"00", x"01", x"03", x"0F", x"0F", x"DF", x"FF", x"FF", x"FF", x"28", x"12", x"08", x"02", x"20", x"00", x"00", x"08", x"80", x"E0", x"F0", x"FD", x"FF", x"FF", x"FF", x"FF", x"40", x"02", x"11", x"40", x"24", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"C8", x"FC", x"FE", x"FF", x"00", x"48", x"00", x"09", x"50", x"80", x"00", x"08", x"01", x"03", x"07", x"07", x"0F", x"1F", x"7F", x"FF", x"10", x"40", x"22", x"08", x"01", x"02", x"40", x"09", x"80", x"80", x"C0", x"E0", x"F8", x"FC", x"FC", x"FE", 
															x"15", x"FD", x"22", x"00", x"08", x"10", x"02", x"40", x"FF", x"68", x"00", x"00", x"00", x"00", x"00", x"00", x"81", x"12", x"6E", x"18", x"04", x"08", x"40", x"00", x"FF", x"7E", x"2C", x"08", x"00", x"00", x"00", x"00", x"42", x"50", x"0E", x"21", x"81", x"04", x"00", x"20", x"FF", x"3F", x"0B", x"01", x"00", x"00", x"00", x"00", x"00", x"81", x"06", x"20", x"72", x"0C", x"42", x"05", x"FF", x"FF", x"FF", x"FF", x"DF", x"07", x"03", x"01", x"01", x"24", x"08", x"03", x"C6", x"18", x"29", x"D0", x"FF", x"FF", x"FF", x"FF", x"FC", x"F0", x"E8", x"C0", x"05", x"43", x"2C", x"F8", x"44", x"01", x"10", x"08", x"FF", x"FE", x"FC", x"50", x"00", x"00", x"00", x"00", x"90", x"B3", x"08", x"50", x"1A", x"04", x"22", x"85", x"FF", x"2F", x"0F", x"1F", x"0F", x"07", x"01", x"00", x"83", x"2C", x"1A", x"4C", x"19", x"B8", x"62", x"90", x"FF", x"FC", x"F2", x"F8", x"F0", x"E8", x"E0", x"80", 
															x"10", x"00", x"84", x"02", x"00", x"24", x"00", x"08", x"01", x"03", x"03", x"01", x"03", x"03", x"01", x"00", x"00", x"22", x"08", x"00", x"41", x"08", x"04", x"20", x"01", x"01", x"07", x"0F", x"07", x"07", x"03", x"01", x"10", x"40", x"C4", x"80", x"00", x"68", x"E0", x"82", x"80", x"C0", x"80", x"80", x"C0", x"E0", x"C0", x"80", x"04", x"30", x"B0", x"20", x"68", x"E1", x"C0", x"88", x"80", x"E0", x"F0", x"E0", x"E0", x"C0", x"80", x"80", x"FF", x"FB", x"FF", x"BF", x"FF", x"EF", x"C5", x"80", x"00", x"04", x"00", x"40", x"00", x"10", x"3A", x"7F", x"FB", x"FF", x"FF", x"E7", x"C3", x"E3", x"87", x"11", x"04", x"00", x"00", x"18", x"3C", x"1C", x"78", x"FE", x"FE", x"BC", x"F8", x"F8", x"F2", x"FC", x"C8", x"04", x"01", x"43", x"07", x"07", x"0F", x"03", x"37", x"FF", x"7F", x"1F", x"1D", x"3F", x"0F", x"87", x"05", x"20", x"80", x"E0", x"E2", x"C0", x"F0", x"F8", x"FE", x"FF", 
															x"FE", x"EE", x"FC", x"FE", x"FC", x"DC", x"FE", x"FF", x"01", x"11", x"03", x"01", x"03", x"23", x"01", x"00", x"FE", x"FC", x"B8", x"F2", x"F0", x"FC", x"F9", x"FE", x"01", x"03", x"47", x"0F", x"0F", x"03", x"07", x"01", x"21", x"87", x"ED", x"FF", x"B6", x"F3", x"E7", x"FD", x"FE", x"7E", x"1B", x"A0", x"49", x"1C", x"1C", x"42", x"01", x"C7", x"9F", x"C5", x"93", x"EF", x"B7", x"F3", x"FE", x"7C", x"71", x"3A", x"7C", x"12", x"48", x"0E", x"00", x"C8", x"B0", x"E2", x"F0", x"BC", x"3A", x"3E", x"FF", x"3F", x"4F", x"1F", x"0F", x"53", x"C5", x"C3", x"01", x"22", x"53", x"3D", x"1F", x"56", x"27", x"73", x"FE", x"FD", x"EC", x"CA", x"F0", x"EB", x"DC", x"8C", x"75", x"3C", x"7F", x"2F", x"17", x"3D", x"39", x"7F", x"8A", x"C3", x"88", x"F0", x"E8", x"C3", x"D6", x"80", x"7F", x"1F", x"4D", x"0F", x"1F", x"8F", x"3F", x"77", x"80", x"E0", x"F2", x"F8", x"E0", x"F2", x"D0", x"C8", 
															x"09", x"FF", x"FF", x"FF", x"DF", x"FF", x"F7", x"FF", x"FF", x"36", x"00", x"00", x"20", x"00", x"08", x"00", x"C9", x"B3", x"EF", x"FF", x"FF", x"FB", x"FF", x"EF", x"FF", x"7E", x"3C", x"10", x"00", x"04", x"00", x"10", x"48", x"DA", x"FE", x"FF", x"DF", x"FF", x"FB", x"FF", x"FF", x"37", x"07", x"01", x"20", x"00", x"04", x"00", x"0A", x"90", x"64", x"08", x"59", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"23", x"01", x"00", x"22", x"09", x"B4", x"C2", x"4F", x"3F", x"9F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FD", x"F8", x"F0", x"C0", x"9B", x"67", x"3F", x"FF", x"FF", x"FB", x"7F", x"FF", x"FF", x"FE", x"FC", x"D0", x"00", x"04", x"80", x"00", x"53", x"C6", x"E8", x"FE", x"F8", x"FD", x"DE", x"FF", x"FF", x"3F", x"1F", x"07", x"0F", x"07", x"23", x"01", x"25", x"57", x"DF", x"3F", x"BE", x"7F", x"BB", x"FF", x"FF", x"FE", x"EC", x"E0", x"E1", x"C0", x"E4", x"80", 
															x"7F", x"37", x"7F", x"FD", x"7F", x"7F", x"FF", x"EF", x"80", x"C8", x"C0", x"82", x"C0", x"C0", x"80", x"10", x"7F", x"7F", x"3D", x"4F", x"BF", x"7F", x"7B", x"FF", x"80", x"C0", x"E2", x"F0", x"E0", x"F0", x"C4", x"80", x"66", x"77", x"F7", x"F3", x"FC", x"7E", x"0E", x"06", x"99", x"99", x"19", x"1F", x"13", x"F3", x"F3", x"FF", x"00", x"70", x"70", x"76", x"67", x"67", x"63", x"00", x"FF", x"8F", x"8F", x"89", x"99", x"99", x"9F", x"FF", x"00", x"18", x"1C", x"1C", x"1C", x"0C", x"00", x"00", x"FF", x"E7", x"E7", x"E7", x"E7", x"FF", x"FF", x"FF", x"00", x"7C", x"7E", x"3E", x"C0", x"E6", x"E6", x"60", x"FF", x"83", x"83", x"FF", x"3F", x"39", x"39", x"FF", x"70", x"7B", x"7B", x"70", x"76", x"77", x"7B", x"38", x"8F", x"8C", x"9C", x"9F", x"99", x"89", x"8F", x"FF", x"E0", x"E6", x"E6", x"E6", x"00", x"3C", x"3C", x"00", x"1F", x"19", x"19", x"19", x"FF", x"C3", x"C3", x"FF", 
															x"40", x"00", x"08", x"00", x"00", x"80", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"C1", x"07", x"04", x"02", x"02", x"04", x"04", x"FF", x"FF", x"3F", x"3C", x"3E", x"3E", x"3C", x"3C", x"01", x"19", x"19", x"11", x"19", x"1A", x"04", x"3C", x"3F", x"27", x"27", x"2F", x"27", x"26", x"3C", x"3C", x"FF", x"FD", x"FF", x"DF", x"FF", x"FF", x"F7", x"FF", x"00", x"02", x"00", x"20", x"00", x"00", x"08", x"00", x"FE", x"D7", x"E3", x"C7", x"AF", x"FE", x"BC", x"FF", x"01", x"28", x"1C", x"3C", x"78", x"19", x"43", x"00", x"FE", x"CF", x"EF", x"C7", x"8F", x"9D", x"FF", x"F7", x"01", x"30", x"10", x"38", x"70", x"62", x"00", x"08", x"4A", x"04", x"90", x"68", x"4C", x"58", x"21", x"03", x"F7", x"FF", x"FF", x"9F", x"BF", x"FF", x"FF", x"FF", 
															x"08", x"10", x"B1", x"40", x"04", x"08", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"4A", x"24", x"8C", x"D1", x"03", x"24", x"18", x"DF", x"BF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"FF", x"FF", x"F7", x"FF", x"FF", x"00", x"00", x"20", x"00", x"00", x"08", x"00", x"00", x"18", x"21", x"2E", x"1F", x"27", x"C2", x"80", x"19", x"FF", x"FE", x"F3", x"FC", x"FD", x"FF", x"FF", x"E6", x"20", x"10", x"C0", x"E0", x"00", x"6D", x"31", x"FC", x"FF", x"FF", x"3F", x"FF", x"FF", x"DF", x"CF", x"57", x"3B", x"FF", x"18", x"66", x"09", x"10", x"00", x"00", x"F4", x"E3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"64", x"00", x"70", x"2C", x"82", x"60", x"40", x"DF", x"FF", x"FF", x"9F", x"DF", x"FF", x"FF", x"FF", x"18", x"85", x"6A", x"42", x"AD", x"19", x"42", x"35", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"03", x"06", x"0A", x"0A", x"18", x"00", x"30", x"20", x"01", x"05", x"05", x"05", x"17", x"1F", x"3F", x"3F", x"80", x"C0", x"A0", x"A0", x"30", x"00", x"18", x"08", x"00", x"40", x"40", x"40", x"D0", x"F0", x"F8", x"F8", x"10", x"22", x"5A", x"2A", x"5A", x"20", x"50", x"20", x"3F", x"3D", x"75", x"75", x"75", x"7F", x"7F", x"7F", x"10", x"88", x"B4", x"A8", x"B4", x"08", x"14", x"08", x"F8", x"78", x"5C", x"5C", x"5C", x"FC", x"FC", x"FC", x"50", x"20", x"50", x"20", x"50", x"21", x"53", x"23", x"7F", x"7F", x"7F", x"7F", x"7F", x"7E", x"7C", x"7C", x"14", x"08", x"14", x"08", x"14", x"08", x"94", x"A8", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"7C", x"7C", x"D1", x"29", x"D1", x"08", x"28", x"10", x"A8", x"50", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"29", x"D1", x"08", x"28", x"10", x"A8", x"50", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"50", x"A0", x"50", x"A0", x"50", x"A0", x"50", x"A0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"15", x"32", x"1D", x"2A", x"1D", x"2E", x"15", x"2E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"50", x"A0", x"51", x"A3", x"53", x"A1", x"51", x"A1", x"FF", x"FF", x"FE", x"FC", x"FC", x"FE", x"FE", x"FE", x"15", x"2E", x"17", x"AF", x"97", x"2B", x"17", x"2B", x"FF", x"FF", x"FF", x"7F", x"7F", x"FF", x"FF", x"FF", x"50", x"A0", x"50", x"A0", x"50", x"20", x"50", x"20", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"14", x"2A", x"14", x"0A", x"14", x"08", x"14", x"08", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"FC", x"FC", x"50", x"20", x"50", x"20", x"50", x"28", x"30", x"E8", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"1F", x"1F", x"14", x"08", x"14", x"08", x"14", x"28", x"18", x"2E", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"F0", x"F0", 
															x"30", x"28", x"11", x"2B", x"13", x"29", x"15", x"09", x"1F", x"1F", x"3E", x"3C", x"3C", x"3E", x"3E", x"1E", x"18", x"28", x"10", x"A8", x"90", x"28", x"50", x"20", x"F0", x"F0", x"F8", x"78", x"78", x"F8", x"F8", x"F0", x"14", x"08", x"14", x"08", x"14", x"08", x"14", x"0A", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"50", x"20", x"50", x"20", x"50", x"20", x"50", x"A0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"15", x"0A", x"54", x"AA", x"54", x"0A", x"04", x"0A", x"1F", x"1F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"50", x"A0", x"54", x"AA", x"D5", x"A0", x"C0", x"E0", x"F0", x"F0", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"54", x"AA", x"54", x"AB", x"0A", x"05", x"07", x"04", x"FF", x"FF", x"FF", x"FF", x"0F", x"0A", x"02", x"00", x"F5", x"FA", x"FD", x"7E", x"A0", x"40", x"C0", x"40", x"FF", x"FF", x"FF", x"FF", x"E0", x"A0", x"80", x"00", 
															x"AA", x"05", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"15", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"55", x"0A", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"0F", x"00", x"00", x"00", x"00", x"00", x"AA", x"55", x"A0", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"F0", x"00", x"00", x"00", x"00", x"00", x"AA", x"55", x"AA", x"55", x"0A", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"00", x"00", x"00", x"AA", x"55", x"AA", x"55", x"A0", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"00", x"00", x"00", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"0A", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"00", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"A0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", 
															x"55", x"0A", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"1F", x"03", x"00", x"00", x"00", x"00", x"00", x"55", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"F0", x"80", x"00", x"00", x"00", x"00", x"00", x"55", x"AA", x"55", x"2A", x"1F", x"06", x"03", x"01", x"FF", x"FF", x"FF", x"7F", x"1F", x"07", x"03", x"01", x"55", x"AA", x"55", x"A8", x"D0", x"C0", x"80", x"00", x"FF", x"FF", x"FF", x"FC", x"F0", x"C0", x"80", x"00", x"00", x"50", x"AA", x"04", x"28", x"40", x"80", x"00", x"00", x"F8", x"FE", x"FC", x"F8", x"E0", x"80", x"00", x"02", x"55", x"AA", x"00", x"00", x"00", x"AA", x"05", x"07", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"80", x"55", x"AA", x"00", x"00", x"01", x"0A", x"A0", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"00", x"00", x"00", x"00", x"01", x"0A", x"00", x"80", x"00", x"00", x"00", x"00", x"03", x"1F", x"7F", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"A0", x"04", x"02", x"00", x"00", x"00", x"00", x"80", x"F0", x"FC", x"FE", x"00", x"00", x"00", x"0A", x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"A0", x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"FF", x"FF", x"FF", x"FF", x"55", x"2A", x"15", x"02", x"00", x"00", x"00", x"00", x"FF", x"7F", x"1F", x"03", x"00", x"00", x"00", x"00", x"54", x"A8", x"50", x"80", x"00", x"00", x"00", x"00", x"FE", x"FC", x"F0", x"80", x"00", x"00", x"00", x"00", x"51", x"AA", x"55", x"AA", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"10", x"28", x"00", x"00", x"00", x"00", x"10", x"10", x"10", x"38", x"54", x"8A", x"44", x"8A", x"44", x"8A", x"44", x"8A", x"7C", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", 
															x"C0", x"00", x"00", x"03", x"0F", x"3F", x"FF", x"F3", x"3F", x"7F", x"FF", x"FC", x"F0", x"C3", x"0C", x"30", x"0F", x"3C", x"F0", x"F0", x"C0", x"00", x"FF", x"FF", x"F0", x"C0", x"00", x"30", x"C0", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"F0", x"C0", x"FF", x"FF", x"FF", x"C3", x"03", x"FF", x"FF", x"00", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"3F", x"FF", x"FF", x"FF", x"DF", x"3F", x"8B", x"87", x"03", x"02", x"81", x"4D", x"3F", x"C7", x"F7", x"79", x"FD", x"FD", x"7E", x"FE", x"86", x"45", x"A6", x"4D", x"2A", x"0C", x"AA", x"55", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AA", x"55", x"AA", x"00", x"00", x"00", x"AA", x"55", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"15", x"AA", x"40", x"2A", x"05", x"00", x"00", x"00", x"3F", x"FF", x"7F", x"3F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"3E", x"3E", x"3E", x"38", x"00", x"FF", x"C7", x"FF", x"C1", x"C1", x"C7", x"FF", x"FF", x"FF", x"FF", x"00", x"30", x"38", x"38", x"18", x"00", x"FF", x"1D", x"FF", x"CF", x"CF", x"CF", x"FF", x"FF", x"FF", x"1D", x"01", x"21", x"61", x"61", x"01", x"01", x"01", x"01", x"FF", x"DF", x"9F", x"9F", x"FF", x"FF", x"FF", x"FF", x"08", x"B2", x"11", x"24", x"01", x"64", x"88", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"61", x"C4", x"24", x"03", x"4A", x"14", x"80", x"32", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"01", x"03", x"07", x"0E", x"1C", x"3C", x"7C", x"00", x"00", x"00", x"00", x"01", x"13", x"33", x"73", x"FF", x"FF", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FD", x"FD", x"FF", x"FF", x"FF", x"6F", x"4F", x"F3", x"F2", x"F2", x"F0", x"F9", x"FB", x"6F", x"4F", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", 
															x"0F", x"0F", x"0F", x"0F", x"0C", x"0C", x"FC", x"FC", x"0F", x"0F", x"00", x"00", x"03", x"03", x"F3", x"F3", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"30", x"30", x"3F", x"3F", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F3", x"F3", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"FF", x"FF", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"80", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FC", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FC", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"03", 
															x"F0", x"F8", x"1C", x"0E", x"07", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FE", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F1", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"FC", x"FC", x"FC", x"E0", x"E0", x"E0", x"FF", x"FF", x"FC", x"0C", x"0C", x"0C", x"FC", x"FC", x"00", x"00", x"03", x"F3", x"F3", x"F3", x"03", x"03", x"FF", x"FF", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF", x"7F", x"3F", x"1F", x"0F", x"F8", x"FC", x"FE", x"FF", x"7F", x"3F", x"10", x"00", x"00", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FF", x"FF", x"03", x"03", x"F3", x"F3", x"F3", x"F3", 
															x"0C", x"0C", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"03", x"03", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"00", x"00", x"F3", x"F3", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"07", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"0E", x"1C", x"F8", x"F0", x"E0", x"C0", x"80", x"00", x"F0", x"E0", x"00", x"00", x"E0", x"C0", x"80", x"00", x"07", x"07", x"0C", x"08", x"38", x"70", x"70", x"E0", x"00", x"00", x"00", x"00", x"27", x"6F", x"4F", x"DF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"BF", x"3F", x"00", x"01", x"01", x"03", x"03", x"07", x"07", x"0E", x"00", x"01", x"01", x"03", x"02", x"06", x"04", x"0D", 
															x"E0", x"C1", x"C1", x"83", x"82", x"06", x"04", x"0C", x"9F", x"BE", x"3E", x"7C", x"7D", x"F9", x"FB", x"F3", x"0E", x"1C", x"1C", x"3C", x"3C", x"7C", x"7C", x"FC", x"09", x"1B", x"13", x"33", x"33", x"73", x"73", x"F3", x"08", x"18", x"1F", x"1F", x"00", x"00", x"00", x"00", x"E7", x"E7", x"C0", x"C0", x"8F", x"8F", x"0F", x"FF", x"30", x"30", x"30", x"3F", x"3F", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"F0", x"F0", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"0C", x"0C", x"00", x"00", x"FF", x"FF", x"F0", x"00", x"03", x"03", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"3F", x"3F", x"30", x"30", x"3F", x"3F", x"03", x"03", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"F0", 
															x"0F", x"0F", x"0C", x"0C", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"00", x"00", x"F3", x"F3", x"F3", x"F3", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"F3", x"F3", x"F3", x"F3", x"F0", x"F0", x"FF", x"FF", x"03", x"03", x"03", x"03", x"FF", x"FF", x"F0", x"F0", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"F0", x"F0", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"7C", x"F0", x"03", x"03", x"F3", x"F3", x"F3", x"F3", x"43", x"0F", x"00", x"00", x"00", x"00", x"03", x"0F", x"0C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"33", x"03", x"0F", x"3C", x"F0", x"C0", x"00", x"00", x"03", x"00", x"00", x"00", x"03", x"0F", x"3F", x"FF", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
	
	constant DONKEY_KONG_JR_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"05", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"00", x"00", x"01", x"C0", x"84", x"A2", x"20", x"1C", x"1F", x"3F", x"7E", x"FF", x"FF", x"FF", x"39", x"1C", x"00", x"00", x"0F", x"1E", x"C7", x"EF", x"3C", x"3C", x"00", x"1F", x"7F", x"FE", x"FE", x"FF", x"FF", x"FF", x"1F", x"71", x"FF", x"0E", x"04", x"00", x"00", x"4E", x"FF", x"8E", x"06", x"F0", x"F8", x"F8", x"F8", x"7E", x"00", x"00", x"00", x"80", x"80", x"F0", x"F0", x"20", x"40", x"80", x"00", x"80", x"E0", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"34", x"1C", x"38", x"E0", x"F0", x"F0", x"F8", x"7C", x"3C", x"1C", x"38", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"08", x"08", x"18", x"00", x"00", x"01", x"03", x"07", x"07", x"07", x"07", x"3C", x"3E", x"42", x"00", x"00", x"00", x"00", x"27", x"03", x"01", x"3D", x"7F", x"7F", x"1F", x"3E", x"3F", x"00", x"1E", x"3D", x"8F", x"DF", x"7F", x"38", x"3F", x"3F", x"FE", x"FD", x"FD", x"FF", x"FF", x"FF", x"FF", x"12", x"1A", x"0C", x"08", x"80", x"88", x"28", x"70", x"ED", x"E5", x"F3", x"F5", x"7E", x"3E", x"3C", x"7E", x"00", x"00", x"00", x"00", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"18", x"0F", x"00", x"00", x"01", x"07", x"0F", x"1F", x"1E", x"0F", x"00", x"00", x"00", x"01", x"09", x"10", x"10", x"30", x"00", x"00", x"00", x"07", x"07", x"0F", x"0F", x"0F", x"78", x"7C", x"1E", x"07", x"07", x"0F", x"20", x"61", x"07", x"03", x"E1", x"F8", x"F8", x"F0", x"39", x"71", x"00", x"1E", x"3D", x"8F", x"DF", x"7F", x"78", x"37", x"3F", x"FE", x"FD", x"FD", x"FF", x"FF", x"FF", x"FF", x"18", x"04", x"00", x"80", x"E0", x"03", x"00", x"9D", x"E6", x"F8", x"FC", x"7F", x"1F", x"FB", x"F0", x"FD", x"00", x"00", x"00", x"00", x"E0", x"E0", x"40", x"80", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"80", x"00", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"80", 
															x"00", x"00", x"00", x"00", x"00", x"38", x"7D", x"68", x"00", x"00", x"00", x"03", x"0F", x"3F", x"7F", x"7F", x"34", x"0E", x"0F", x"2B", x"40", x"80", x"E0", x"00", x"33", x"01", x"00", x"34", x"7F", x"FF", x"EF", x"00", x"00", x"00", x"01", x"03", x"31", x"3B", x"1F", x"1F", x"00", x"03", x"0F", x"9F", x"FF", x"FF", x"EF", x"EF", x"1F", x"3B", x"F8", x"FD", x"FF", x"3C", x"00", x"00", x"E7", x"C7", x"07", x"02", x"00", x"C3", x"80", x"00", x"03", x"05", x"E6", x"B3", x"F9", x"FC", x"8C", x"1C", x"03", x"E7", x"F7", x"B7", x"BF", x"FF", x"FF", x"FF", x"18", x"E0", x"40", x"C8", x"1C", x"3C", x"70", x"00", x"FE", x"F8", x"80", x"38", x"FC", x"FC", x"F0", x"00", x"40", x"C0", x"60", x"C0", x"80", x"00", x"00", x"00", x"40", x"C0", x"E0", x"C0", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"0C", x"1E", x"1F", x"1E", x"0C", x"00", x"00", x"0F", x"1F", x"1F", x"1F", x"1F", x"0D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"02", x"03", x"03", x"01", x"01", x"C7", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"01", x"01", x"01", x"0B", x"04", x"00", x"00", x"01", x"3E", x"1E", x"1E", x"04", x"03", x"02", x"01", x"01", x"00", x"7C", x"FC", x"68", x"F4", x"FE", x"86", x"8F", x"F8", x"FD", x"E3", x"C3", x"EB", x"FF", x"FF", x"FE", x"FD", x"E3", x"FF", x"0E", x"06", x"04", x"01", x"38", x"FE", x"1C", x"00", x"F1", x"79", x"FB", x"F1", x"F8", x"00", x"00", x"00", x"00", x"38", x"78", x"20", x"00", x"00", x"C0", x"F0", x"D0", x"F8", x"F8", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"E0", x"F0", x"00", 
															x"00", x"01", x"0B", x"0E", x"06", x"19", x"17", x"1F", x"03", x"07", x"0E", x"0C", x"0F", x"1F", x"3F", x"3F", x"0F", x"00", x"10", x"1E", x"0F", x"07", x"03", x"00", x"3F", x"1F", x"0F", x"01", x"00", x"00", x"00", x"00", x"00", x"C0", x"EB", x"BB", x"31", x"CC", x"F4", x"FD", x"E0", x"F0", x"3B", x"1F", x"FF", x"FF", x"FC", x"FD", x"F9", x"00", x"00", x"02", x"CC", x"C0", x"E0", x"E0", x"FB", x"FF", x"FF", x"FF", x"3F", x"3F", x"1E", x"00", x"00", x"00", x"C0", x"40", x"C0", x"00", x"00", x"E0", x"00", x"00", x"C0", x"C0", x"C0", x"00", x"00", x"E0", x"60", x"E0", x"00", x"00", x"08", x"08", x"08", x"10", x"E0", x"E0", x"00", x"80", x"D8", x"F8", x"F8", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"01", x"0B", x"0E", x"06", x"19", x"17", x"1F", x"03", x"07", x"0E", x"0C", x"0F", x"1F", x"3F", x"3F", x"0F", x"00", x"10", x"1E", x"0F", x"07", x"03", x"00", x"3F", x"1F", x"0F", x"01", x"00", x"00", x"00", x"00", x"03", x"C3", x"EA", x"BB", x"30", x"CD", x"F5", x"FC", x"E3", x"F3", x"3F", x"1F", x"FE", x"FD", x"FD", x"FF", x"F8", x"01", x"02", x"08", x"C0", x"C0", x"E0", x"E0", x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"1B", x"03", x"C0", x"40", x"C0", x"80", x"00", x"E0", x"60", x"E0", x"C0", x"C0", x"C0", x"80", x"00", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"C0", x"80", x"00", x"80", x"C0", x"C0", x"80", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"74", x"64", x"70", x"20", x"00", x"00", x"00", x"00", x"74", x"66", x"77", x"27", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"03", x"01", x"00", x"00", x"00", x"01", x"03", x"03", x"03", x"01", x"00", x"01", x"0C", x"1F", x"17", x"18", x"3C", x"36", x"00", x"00", x"0F", x"DF", x"FF", x"EF", x"CF", x"CF", x"3B", x"3C", x"1B", x"1C", x"0D", x"07", x"00", x"C0", x"47", x"03", x"64", x"E3", x"F2", x"F8", x"E0", x"C0", x"C0", x"70", x"B8", x"F4", x"FE", x"7C", x"3C", x"78", x"78", x"7C", x"2C", x"9C", x"FC", x"FB", x"FB", x"F7", x"F0", x"60", x"F4", x"F8", x"E0", x"C0", x"01", x"00", x"EF", x"9F", x"08", x"07", x"1F", x"3F", x"03", x"00", x"00", x"00", x"00", x"0E", x"26", x"2E", x"04", x"00", x"00", x"00", x"00", x"0E", x"26", x"6E", x"E4", x"E0", x"00", x"00", x"00", x"00", x"30", x"F0", x"80", x"00", x"E0", x"C0", x"00", x"30", x"F0", x"F0", x"80", x"00", 
															x"00", x"00", x"00", x"00", x"58", x"E8", x"D8", x"70", x"00", x"00", x"00", x"00", x"58", x"FF", x"FF", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"3A", x"3E", x"1E", x"33", x"20", x"27", x"03", x"01", x"05", x"01", x"01", x"FC", x"FF", x"FF", x"1F", x"00", x"0F", x"0C", x"0F", x"04", x"1B", x"F0", x"FF", x"7F", x"30", x"13", x"70", x"FB", x"7C", x"F0", x"00", x"70", x"50", x"70", x"38", x"CC", x"04", x"E4", x"C0", x"80", x"A0", x"80", x"F8", x"3F", x"FF", x"FF", x"F8", x"00", x"F0", x"30", x"70", x"E0", x"C0", x"0F", x"FF", x"FE", x"08", x"C8", x"8E", x"1F", x"3E", x"0F", x"00", x"00", x"00", x"00", x"00", x"08", x"0E", x"1F", x"00", x"00", x"00", x"00", x"00", x"F8", x"FE", x"FF", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"0B", x"1D", x"1B", x"0E", x"00", x"00", x"00", x"00", x"0B", x"1F", x"1F", x"0F", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"04", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"05", x"07", x"03", x"01", x"00", x"00", x"0E", x"0A", x"0E", x"1E", x"33", x"20", x"20", x"03", x"01", x"C5", x"E1", x"FF", x"FC", x"FF", x"7F", x"27", x"18", x"07", x"0C", x"0F", x"04", x"83", x"00", x"3F", x"3F", x"D8", x"F3", x"F0", x"FB", x"8C", x"00", x"70", x"F8", x"B8", x"F8", x"78", x"8C", x"04", x"04", x"80", x"00", x"40", x"01", x"8F", x"7F", x"FF", x"FF", x"E4", x"18", x"E0", x"30", x"70", x"E5", x"C7", x"00", x"FE", x"FC", x"1F", x"CF", x"8F", x"1F", x"27", x"00", x"00", x"60", x"5C", x"6C", x"38", x"00", x"00", x"00", x"00", x"60", x"7C", x"FC", x"F8", x"E0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"0B", x"0F", x"07", x"03", x"03", x"07", x"07", x"07", x"0F", x"0F", x"07", x"03", x"00", x"01", x"0B", x"2E", x"26", x"3F", x"37", x"38", x"03", x"07", x"1E", x"1C", x"5F", x"DF", x"DF", x"DF", x"1F", x"0C", x"1F", x"3E", x"1F", x"06", x"03", x"00", x"EF", x"F3", x"A0", x"01", x"00", x"39", x"1C", x"3E", x"00", x"C0", x"E8", x"BA", x"32", x"6E", x"76", x"0E", x"E0", x"F0", x"3C", x"1C", x"FD", x"FD", x"FD", x"FD", x"FC", x"18", x"FC", x"1E", x"BC", x"70", x"E0", x"00", x"FB", x"E7", x"02", x"E0", x"40", x"8E", x"1C", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"00", x"00", x"00", x"00", x"68", x"F8", x"70", x"60", x"E0", x"F0", x"F0", x"70", x"78", x"F8", x"70", x"60", 
															x"06", x"0F", x"05", x"07", x"87", x"4E", x"57", x"23", x"02", x"01", x"01", x"07", x"83", x"4C", x"57", x"23", x"3C", x"7C", x"F8", x"E0", x"80", x"2A", x"FE", x"FC", x"3C", x"78", x"E0", x"80", x"00", x"00", x"AA", x"FC", x"00", x"01", x"01", x"03", x"87", x"4F", x"37", x"03", x"00", x"00", x"00", x"02", x"83", x"4D", x"37", x"03", x"80", x"C0", x"40", x"FC", x"FE", x"FE", x"FE", x"FC", x"80", x"40", x"40", x"7C", x"FE", x"54", x"AA", x"FC", x"92", x"54", x"38", x"FE", x"38", x"54", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"81", x"81", x"81", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"09", x"01", x"02", x"01", x"09", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"60", x"C3", x"E7", x"C7", x"EF", x"CE", x"DC", x"00", x"40", x"81", x"C3", x"83", x"C7", x"86", x"CC", x"DE", x"FB", x"7F", x"20", x"40", x"80", x"60", x"10", x"DE", x"D9", x"68", x"20", x"40", x"80", x"60", x"10", x"00", x"70", x"F8", x"F8", x"F8", x"F8", x"FE", x"FB", x"00", x"50", x"B8", x"D8", x"B8", x"D8", x"BE", x"D1", x"FE", x"F8", x"70", x"20", x"40", x"40", x"20", x"10", x"F0", x"D8", x"60", x"20", x"40", x"40", x"20", x"10", x"00", x"00", x"00", x"00", x"1E", x"3F", x"7D", x"78", x"00", x"00", x"01", x"00", x"00", x"20", x"7C", x"78", x"7C", x"FB", x"FF", x"FF", x"5F", x"1F", x"1F", x"1F", x"7C", x"FE", x"FF", x"FE", x"7C", x"60", x"E0", x"E1", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"7C", x"82", x"01", x"82", x"7C", x"00", x"00", x"00", x"00", x"21", x"A2", x"A3", x"B3", x"8F", x"27", x"FE", x"10", x"19", x"5A", x"DF", x"4F", x"73", x"DB", x"02", 
															x"00", x"00", x"00", x"01", x"03", x"0F", x"BF", x"FF", x"00", x"00", x"00", x"00", x"00", x"0C", x"BE", x"FF", x"FF", x"FF", x"7F", x"3F", x"7F", x"F8", x"00", x"00", x"F3", x"FF", x"63", x"FE", x"0D", x"F8", x"00", x"00", x"00", x"00", x"00", x"80", x"70", x"60", x"D0", x"C0", x"00", x"00", x"00", x"00", x"30", x"38", x"7C", x"FE", x"C0", x"C0", x"E0", x"F0", x"E0", x"00", x"00", x"00", x"FF", x"F0", x"7E", x"F8", x"E0", x"00", x"00", x"00", x"00", x"78", x"FC", x"7E", x"7F", x"3F", x"3F", x"9F", x"00", x"78", x"FC", x"0E", x"7E", x"3C", x"0C", x"9E", x"FF", x"FF", x"FF", x"0F", x"1F", x"0F", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"5F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"70", x"60", x"D0", x"00", x"00", x"00", x"00", x"00", x"3F", x"3E", x"7E", x"C0", x"C0", x"C0", x"E0", x"F0", x"80", x"00", x"00", x"FC", x"F8", x"FC", x"FE", x"FF", x"80", x"00", x"00", 
															x"00", x"00", x"03", x"43", x"61", x"77", x"7F", x"7F", x"00", x"00", x"03", x"47", x"43", x"57", x"77", x"74", x"7E", x"3E", x"0E", x"01", x"00", x"00", x"00", x"00", x"7C", x"3C", x"0F", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"E0", x"E1", x"C3", x"F7", x"FF", x"FF", x"00", x"00", x"E0", x"F1", x"E1", x"F5", x"F7", x"97", x"BF", x"BE", x"38", x"40", x"00", x"00", x"00", x"00", x"1F", x"1E", x"F8", x"F0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"03", x"04", x"0B", x"17", x"00", x"00", x"07", x"08", x"93", x"27", x"4C", x"5A", x"17", x"0B", x"04", x"03", x"00", x"00", x"00", x"00", x"5A", x"4C", x"27", x"13", x"08", x"27", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"20", x"D0", x"E0", x"00", x"04", x"E0", x"10", x"C8", x"E4", x"32", x"52", x"E8", x"D0", x"20", x"C0", x"00", x"00", x"00", x"00", x"5A", x"32", x"E4", x"C8", x"12", x"E0", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"03", x"04", x"0A", x"00", x"00", x"00", x"20", x"00", x"00", x"03", x"07", x"0A", x"04", x"03", x"00", x"00", x"00", x"00", x"00", x"07", x"03", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"20", x"50", x"00", x"00", x"00", x"02", x"00", x"00", x"C0", x"E0", x"50", x"20", x"C0", x"00", x"00", x"00", x"00", x"00", x"E0", x"C0", x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"04", x"00", x"00", x"01", x"23", x"04", x"0B", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0D", x"0F", x"4B", x"04", x"0B", x"21", x"02", x"00", x"00", x"11", x"0C", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"C0", x"E2", x"90", x"E8", x"00", x"00", x"00", x"80", x"40", x"60", x"70", x"58", x"F8", x"E8", x"94", x"E0", x"D2", x"00", x"00", x"00", x"44", x"18", x"70", x"60", x"40", x"80", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"05", x"00", x"00", x"00", x"00", x"02", x"01", x"03", x"07", x"05", x"02", x"01", x"00", x"01", x"00", x"00", x"00", x"07", x"03", x"11", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C8", x"20", x"D0", x"00", x"00", x"00", x"00", x"00", x"C8", x"E0", x"70", x"D0", x"20", x"C8", x"00", x"00", x"00", x"00", x"00", x"74", x"E0", x"C8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"F2", x"20", x"04", x"01", x"09", x"00", x"00", x"47", x"FD", x"3F", x"1B", x"1F", x"17", x"1C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"78", x"78", x"BC", x"00", x"00", x"00", x"00", x"30", x"F2", x"FF", x"BF", x"01", x"80", x"E0", x"80", 
															x"00", x"00", x"00", x"00", x"00", x"1C", x"00", x"06", x"00", x"00", x"00", x"00", x"3E", x"63", x"3F", x"19", x"40", x"F2", x"38", x"1F", x"07", x"01", x"00", x"00", x"5F", x"FD", x"3F", x"1F", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"78", x"F8", x"BC", x"00", x"00", x"00", x"00", x"B0", x"F2", x"FF", x"BF", x"01", x"80", x"E0", x"80", x"00", x"01", x"01", x"01", x"03", x"21", x"09", x"01", x"00", x"01", x"41", x"61", x"73", x"5F", x"37", x"3F", x"00", x"01", x"07", x"07", x"02", x"00", x"00", x"00", x"18", x"01", x"07", x"04", x"00", x"01", x"00", x"00", x"00", x"E0", x"C0", x"C0", x"E0", x"C2", x"C8", x"C0", x"00", x"E0", x"C1", x"C3", x"E7", x"FD", x"F6", x"FE", x"80", x"E0", x"F0", x"F0", x"20", x"00", x"00", x"00", x"80", x"E0", x"F0", x"90", x"80", x"C0", x"80", x"00", 
															x"3C", x"7E", x"C3", x"81", x"81", x"C3", x"7E", x"3C", x"3C", x"42", x"81", x"00", x"00", x"81", x"42", x"3C", x"00", x"18", x"3C", x"66", x"66", x"3C", x"18", x"00", x"00", x"18", x"24", x"42", x"42", x"24", x"18", x"00", x"00", x"00", x"00", x"10", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"10", x"28", x"10", x"00", x"00", x"99", x"42", x"00", x"80", x"01", x"00", x"42", x"99", x"08", x"42", x"00", x"80", x"01", x"00", x"42", x"10", x"00", x"00", x"03", x"06", x"0C", x"0C", x"18", x"20", x"FF", x"FF", x"03", x"07", x"0D", x"0D", x"19", x"39", x"20", x"18", x"0C", x"0C", x"06", x"03", x"00", x"00", x"39", x"19", x"0D", x"0D", x"07", x"03", x"FF", x"FF", x"00", x"00", x"C0", x"60", x"30", x"30", x"18", x"04", x"FF", x"FF", x"C0", x"E0", x"B0", x"B0", x"98", x"9C", x"04", x"18", x"30", x"30", x"60", x"C0", x"00", x"00", x"9C", x"98", x"B0", x"B0", x"E0", x"C0", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0E", x"00", x"00", x"00", x"00", x"FF", x"FF", x"03", x"0F", x"38", x"40", x"40", x"38", x"0E", x"03", x"00", x"00", x"39", x"71", x"71", x"39", x"0F", x"03", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"70", x"00", x"00", x"00", x"00", x"FF", x"FF", x"C0", x"F0", x"1C", x"02", x"02", x"1C", x"70", x"C0", x"00", x"00", x"9C", x"8E", x"8E", x"9C", x"F0", x"C0", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"38", x"38", x"0F", x"00", x"00", x"FF", x"FF", x"0F", x"F9", x"F9", x"0F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"1C", x"1C", x"F0", x"00", x"00", x"FF", x"FF", x"F0", x"9F", x"9F", x"F0", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"1F", x"00", x"00", x"0C", x"1E", x"01", x"07", x"0C", x"18", x"1F", x"1F", x"1F", x"0F", x"07", x"03", x"00", x"00", x"19", x"1F", x"1F", x"0F", x"07", x"03", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"E0", x"F0", x"F8", x"00", x"00", x"B0", x"F8", x"C0", x"E0", x"F0", x"F8", x"F8", x"F8", x"F8", x"F0", x"E0", x"C0", x"00", x"00", x"F8", x"F8", x"F8", x"F0", x"E0", x"C0", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E7", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"27", x"FF", x"80", x"1F", x"03", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"3F", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"38", x"F0", x"E0", x"00", x"00", x"00", x"00", x"0C", x"3C", x"FC", x"F8", x"C0", x"0C", x"F8", x"E0", x"00", x"00", x"00", x"00", x"F8", x"FC", x"FE", x"FE", x"FC", x"F0", x"00", x"00", x"00", x"00", x"00", x"0C", x"0E", x"07", x"0F", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"3F", x"7C", x"7C", x"78", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"38", x"70", x"80", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F0", x"F8", x"F8", x"F8", x"78", x"10", x"00", x"00", x"FC", x"FE", x"FE", x"FE", x"7E", x"1C", x"00", x"00", 
															x"7F", x"FF", x"FF", x"EE", x"E4", x"44", x"44", x"40", x"00", x"10", x"21", x"13", x"1B", x"BB", x"00", x"00", x"FE", x"FF", x"FF", x"F7", x"72", x"62", x"22", x"02", x"10", x"08", x"44", x"08", x"8D", x"9D", x"00", x"00", x"18", x"18", x"00", x"10", x"10", x"10", x"10", x"10", x"66", x"66", x"3C", x"18", x"18", x"18", x"18", x"18", x"10", x"10", x"10", x"10", x"00", x"20", x"02", x"04", x"18", x"18", x"18", x"18", x"3C", x"5E", x"7E", x"3C", x"0F", x"1F", x"1E", x"24", x"26", x"70", x"00", x"1F", x"0F", x"1F", x"01", x"1B", x"19", x"0F", x"1F", x"03", x"3F", x"3F", x"7F", x"7E", x"7F", x"3F", x"3C", x"3E", x"00", x"00", x"60", x"7F", x"7F", x"3F", x"04", x"00", x"00", x"E0", x"00", x"80", x"40", x"F0", x"00", x"38", x"00", x"E0", x"80", x"70", x"B8", x"01", x"C3", x"07", x"FC", x"F8", x"E0", x"F4", x"FC", x"F8", x"30", x"00", x"03", x"00", x"20", x"F0", x"F0", x"E0", x"00", x"00", 
															x"00", x"07", x"0F", x"0F", x"12", x"13", x"38", x"00", x"00", x"07", x"0F", x"00", x"0D", x"0C", x"07", x"0F", x"1F", x"1F", x"3F", x"FF", x"FF", x"BF", x"41", x"01", x"10", x"10", x"38", x"7F", x"7F", x"3F", x"00", x"00", x"00", x"80", x"F0", x"00", x"40", x"20", x"78", x"00", x"00", x"80", x"F0", x"C0", x"B8", x"DC", x"81", x"E3", x"F8", x"FC", x"A0", x"E0", x"F0", x"F0", x"C0", x"E0", x"07", x"03", x"E0", x"E0", x"F0", x"F0", x"C0", x"00", x"1E", x"3F", x"3C", x"49", x"4C", x"E1", x"00", x"39", x"1E", x"3F", x"03", x"36", x"33", x"1E", x"3F", x"3F", x"7F", x"7F", x"7D", x"7F", x"3F", x"1E", x"1C", x"1E", x"00", x"00", x"47", x"7F", x"3F", x"1E", x"00", x"00", x"00", x"C0", x"00", x"00", x"80", x"E0", x"00", x"00", x"08", x"C8", x"04", x"E2", x"71", x"02", x"84", x"08", x"E0", x"E0", x"C0", x"E0", x"E0", x"E0", x"F0", x"00", x"1C", x"1C", x"C8", x"E0", x"E0", x"E0", x"00", x"00", 
															x"0F", x"1F", x"1E", x"24", x"26", x"70", x"00", x"1F", x"0F", x"1F", x"01", x"1B", x"19", x"0F", x"1F", x"04", x"3F", x"3F", x"3E", x"FF", x"FC", x"F8", x"40", x"01", x"02", x"03", x"21", x"70", x"7B", x"3B", x"01", x"00", x"00", x"E0", x"00", x"80", x"40", x"F0", x"00", x"80", x"00", x"E0", x"C0", x"70", x"B8", x"00", x"C0", x"00", x"E0", x"E0", x"E0", x"E0", x"60", x"00", x"80", x"E0", x"40", x"38", x"F8", x"E2", x"E2", x"C1", x"F2", x"1C", x"07", x"0F", x"0A", x"10", x"36", x"33", x"01", x"6F", x"07", x"0F", x"15", x"0F", x"09", x"0C", x"07", x"04", x"7F", x"1B", x"0F", x"1F", x"7F", x"7E", x"1C", x"00", x"06", x"0F", x"0F", x"1F", x"0F", x"02", x"00", x"00", x"E0", x"F0", x"50", x"08", x"6C", x"CC", x"80", x"F6", x"E0", x"F0", x"A8", x"F0", x"90", x"30", x"E0", x"20", x"FE", x"D8", x"F3", x"FF", x"FE", x"3E", x"00", x"00", x"60", x"F0", x"F0", x"F8", x"F0", x"30", x"00", x"00", 
															x"00", x"00", x"79", x"F9", x"F3", x"FF", x"7B", x"3F", x"00", x"01", x"00", x"00", x"00", x"1E", x"7F", x"3E", x"3F", x"3F", x"7B", x"7F", x"FB", x"F1", x"79", x"38", x"3C", x"3E", x"7F", x"7E", x"18", x"00", x"00", x"00", x"00", x"00", x"80", x"B0", x"B8", x"C6", x"93", x"F7", x"C0", x"E0", x"40", x"00", x"00", x"3A", x"EF", x"4B", x"E3", x"F7", x"93", x"C6", x"B8", x"B0", x"80", x"00", x"5F", x"4B", x"EF", x"3A", x"00", x"00", x"60", x"C0", x"7B", x"07", x"02", x"00", x"00", x"01", x"01", x"01", x"7B", x"3F", x"7E", x"7C", x"FC", x"FF", x"FF", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"3F", x"0F", x"01", x"00", x"00", x"00", x"00", x"01", x"00", x"9B", x"36", x"BF", x"F1", x"BF", x"9F", x"C0", x"1F", x"BF", x"64", x"E0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"78", x"7F", x"1F", x"01", x"D4", x"FF", x"3F", x"9F", x"07", x"80", x"E0", x"7E", x"FC", 
															x"0E", x"1F", x"83", x"A0", x"E0", x"B0", x"30", x"70", x"0E", x"9F", x"C3", x"E1", x"E1", x"F3", x"FF", x"FF", x"E0", x"C0", x"E0", x"F1", x"FE", x"FC", x"F8", x"01", x"FF", x"BF", x"1F", x"0E", x"01", x"03", x"07", x"01", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"E0", x"F0", x"F0", x"F8", x"F8", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"20", x"70", x"F0", x"E0", x"80", x"00", x"80", x"C0", x"E0", x"F0", x"F0", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"03", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"1F", x"1F", x"1F", x"0F", x"07", x"03", x"00", x"00", x"00", x"00", x"01", x"02", x"04", x"04", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"04", x"00", x"00", x"03", x"07", x"0A", x"00", x"00", x"07", x"03", x"01", x"03", x"07", x"0F", x"00", x"00", 
															x"00", x"00", x"78", x"EC", x"76", x"A0", x"DC", x"F8", x"00", x"00", x"78", x"FC", x"FE", x"FC", x"FC", x"F9", x"10", x"34", x"20", x"40", x"00", x"00", x"00", x"00", x"F3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"82", x"81", x"01", x"02", x"01", x"00", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"4C", x"FA", x"BE", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"0F", x"5F", x"CE", x"00", x"00", x"07", x"0F", x"1F", x"3F", x"7C", x"FC", x"CF", x"7E", x"FF", x"E0", x"DF", x"3F", x"3F", x"0F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"55", x"AA", x"FE", x"EE", x"7D", x"83", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"37", x"0F", x"05", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"1F", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"30", x"78", x"FD", x"B9", x"00", x"00", x"F0", x"F8", x"FC", x"FE", x"9F", x"9F", x"F9", x"3F", x"FF", x"03", x"FD", x"FE", x"FE", x"F8", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"55", x"AA", x"FF", x"EF", x"7C", x"83", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D8", x"E0", x"40", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1B", x"37", x"82", x"00", x"00", x"00", x"00", x"0F", x"1F", x"3F", x"9F", x"9D", x"0F", x"84", x"86", x"82", x"01", x"00", x"00", x"DF", x"CF", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"80", x"08", x"04", x"82", x"01", x"01", x"FF", x"FC", x"F8", x"F8", x"FC", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"65", x"BF", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"C0", x"60", x"F0", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"F0", x"E0", x"00", x"00", x"00", x"80", x"00", x"00", x"F0", x"F8", x"FC", x"FC", x"FE", x"FE", x"FE", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"00", x"80", x"C0", x"A0", x"80", x"80", x"80", x"80", x"00", x"80", x"C0", x"E0", x"00", x"00", x"00", x"06", x"0F", x"5F", x"CE", x"CF", x"00", x"07", x"0F", x"1F", x"3F", x"7C", x"FC", x"FF", x"7E", x"FF", x"F7", x"A2", x"77", x"3F", x"0F", x"00", x"FF", x"CF", x"88", x"DD", x"C8", x"F0", x"FF", x"FF", x"00", x"00", x"00", x"30", x"78", x"FD", x"B9", x"FB", x"00", x"F0", x"F8", x"FC", x"FE", x"9F", x"9F", x"FF", x"3E", x"FF", x"77", x"23", x"76", x"FC", x"F0", x"00", x"FF", x"F3", x"89", x"DD", x"8B", x"0F", x"FF", x"FF", 
															x"70", x"FC", x"FE", x"FE", x"FF", x"7F", x"3E", x"1C", x"00", x"00", x"40", x"40", x"60", x"30", x"1E", x"00", x"02", x"06", x"02", x"02", x"02", x"02", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"09", x"01", x"02", x"04", x"08", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"05", x"09", x"09", x"0F", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"09", x"09", x"06", x"09", x"09", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"26", x"69", x"21", x"22", x"24", x"28", x"2F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"26", x"69", x"28", x"2E", x"29", x"29", x"26", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"22", x"55", x"55", x"55", x"55", x"55", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"78", x"C4", x"E4", x"78", x"86", x"86", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3E", x"60", x"C0", x"DE", x"C6", x"66", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"06", x"06", x"06", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"0E", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"65", x"79", x"65", x"65", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E4", x"96", x"96", x"97", x"96", x"E6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"59", x"59", x"59", x"59", x"D9", x"4E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"70", x"70", x"3C", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"28", x"28", x"28", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"0E", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"28", x"28", x"28", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"70", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"3C", x"38", x"30", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"10", x"10", x"70", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3F", x"7F", x"E0", x"C0", x"C0", x"C0", x"CC", x"CF", x"3F", x"60", x"C1", x"83", x"87", x"87", x"8F", x"8F", x"CF", x"DF", x"DF", x"DF", x"CF", x"C7", x"C3", x"C0", x"8F", x"9F", x"9F", x"9F", x"8F", x"87", x"83", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"81", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"7F", x"3F", x"81", x"81", x"81", x"80", x"83", x"C7", x"60", x"3F", x"FF", x"FF", x"11", x"89", x"5D", x"21", x"01", x"E3", x"FF", x"00", x"FC", x"FE", x"FC", x"FC", x"F8", x"F2", x"CB", x"DF", x"9F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"3F", x"1F", x"0F", x"1F", x"3F", x"7F", x"7F", x"FF", x"3E", x"1E", x"1E", x"3E", x"7E", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"59", x"03", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"FF", 
															x"FF", x"FF", x"8F", x"99", x"B0", x"A3", x"B2", x"B0", x"FF", x"00", x"0F", x"1F", x"3F", x"7C", x"7C", x"7F", x"81", x"B0", x"FF", x"FF", x"BF", x"C7", x"F0", x"FF", x"7F", x"4F", x"08", x"5D", x"48", x"78", x"7F", x"7F", x"D5", x"AA", x"80", x"88", x"C1", x"BE", x"90", x"E4", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"F8", x"FD", x"C0", x"80", x"80", x"80", x"FF", x"FF", x"7F", x"7F", x"40", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"F9", x"CD", x"87", x"63", x"27", x"07", x"FF", x"00", x"F8", x"FC", x"FE", x"9E", x"9E", x"FE", x"C1", x"07", x"FF", x"FF", x"FF", x"F9", x"03", x"FF", x"FE", x"F8", x"88", x"DC", x"88", x"06", x"FE", x"FE", x"55", x"AB", x"81", x"89", x"41", x"3F", x"05", x"13", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"0F", x"5F", x"03", x"01", x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"02", x"00", x"00", x"00", x"00", x"FF", 
															x"FF", x"FF", x"88", x"91", x"BA", x"84", x"80", x"C6", x"FF", x"00", x"3F", x"7F", x"3F", x"3F", x"1F", x"4F", x"D3", x"FB", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FC", x"F8", x"F0", x"F8", x"FC", x"FE", x"FE", x"FF", x"7C", x"78", x"78", x"7C", x"7E", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"9A", x"C0", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"FF", x"FC", x"FE", x"07", x"03", x"03", x"03", x"33", x"F3", x"FC", x"06", x"83", x"C1", x"E1", x"E1", x"F1", x"F1", x"F3", x"FB", x"FB", x"FB", x"F3", x"E3", x"C3", x"03", x"F1", x"F9", x"F9", x"F9", x"F1", x"E1", x"C1", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"03", x"03", x"03", x"03", x"07", x"FE", x"FC", x"81", x"81", x"81", x"01", x"C1", x"E3", x"06", x"FC", 
															x"0F", x"1F", x"1E", x"24", x"26", x"70", x"00", x"1F", x"0F", x"1F", x"01", x"1B", x"19", x"0F", x"1F", x"04", x"3F", x"3F", x"3E", x"FF", x"FC", x"F8", x"40", x"01", x"02", x"03", x"21", x"70", x"7B", x"3B", x"01", x"00", x"00", x"E0", x"00", x"80", x"40", x"F0", x"00", x"80", x"00", x"E0", x"80", x"70", x"B8", x"00", x"C0", x"00", x"E0", x"E0", x"E0", x"E0", x"60", x"00", x"80", x"E0", x"40", x"38", x"F8", x"E2", x"E2", x"C1", x"E2", x"1C", x"3F", x"60", x"5F", x"5E", x"5D", x"5C", x"5E", x"5E", x"00", x"1F", x"20", x"21", x"22", x"23", x"21", x"21", x"5E", x"5E", x"5E", x"2E", x"13", x"0C", x"03", x"03", x"21", x"21", x"21", x"11", x"0C", x"03", x"00", x"00", x"FC", x"06", x"FA", x"7A", x"BA", x"3A", x"7A", x"7A", x"00", x"F8", x"04", x"84", x"44", x"C4", x"84", x"84", x"7A", x"3A", x"7A", x"34", x"C8", x"30", x"C0", x"C0", x"84", x"C4", x"84", x"C8", x"30", x"C0", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"1F", x"00", x"00", x"0C", x"1E", x"01", x"07", x"0C", x"18", x"1F", x"1F", x"1F", x"0F", x"07", x"03", x"00", x"00", x"19", x"1F", x"1F", x"0F", x"07", x"03", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"E0", x"F0", x"F8", x"00", x"00", x"B0", x"F8", x"C0", x"E0", x"F0", x"F8", x"F8", x"F8", x"F8", x"F0", x"E0", x"C0", x"00", x"00", x"F8", x"F8", x"F8", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E7", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"27", x"FF", x"80", x"1F", x"03", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"3F", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"38", x"F0", x"E0", x"00", x"00", x"00", x"00", x"0C", x"3C", x"FC", x"F8", x"C0", x"0C", x"F8", x"E0", x"00", x"00", x"00", x"00", x"F8", x"FC", x"FE", x"FE", x"FC", x"F0", x"00", x"00", 
															x"00", x"00", x"00", x"06", x"07", x"03", x"07", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"3E", x"3E", x"3C", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"1E", x"00", x"00", x"00", x"00", x"10", x"10", x"10", x"14", x"1C", x"38", x"D0", x"60", x"18", x"18", x"18", x"18", x"00", x"00", x"18", x"FC", x"78", x"7C", x"7C", x"7C", x"3C", x"18", x"10", x"10", x"FE", x"FF", x"7F", x"7F", x"3F", x"1E", x"18", x"18", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"10", x"10", x"10", x"10", x"30", x"74", x"76", x"D2", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"FF", x"00", x"30", x"04", x"00", x"00", x"00", x"E1", x"FF", x"FF", x"FF", x"FF", x"FD", x"83", x"FD", x"FF", x"0F", x"3F", x"7F", x"FF", x"FF", x"F7", x"61", x"00", x"00", x"04", x"08", x"10", x"00", x"00", x"08", x"3E", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"EF", x"C6", x"00", x"00", x"00", x"22", x"0C", x"00", x"00", x"10", x"39", x"F0", x"FC", x"FE", x"FF", x"FF", x"EF", x"C6", x"00", x"00", x"30", x"08", x"00", x"00", x"00", x"10", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"BF", x"DB", x"E7", x"FF", x"80", x"C3", x"FF", x"BD", x"CE", x"B3", x"DF", x"FF", x"00", x"00", x"00", x"42", x"31", x"4C", x"20", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"14", x"14", x"08", x"08", x"14", x"14", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"08", x"14", x"14", x"08", x"08", x"1C", x"3E", x"1C", x"00", x"00", x"24", x"00", x"00", x"24", x"00", x"00", x"81", x"81", x"7E", x"24", x"24", x"7E", x"81", x"81", 
															x"7E", x"BF", x"FF", x"2C", x"2C", x"2C", x"2C", x"2C", x"00", x"40", x"00", x"10", x"10", x"10", x"10", x"10", x"FF", x"00", x"FF", x"3C", x"18", x"18", x"18", x"18", x"00", x"FF", x"00", x"C3", x"04", x"04", x"04", x"04", x"18", x"18", x"18", x"18", x"3C", x"FF", x"FF", x"00", x"04", x"04", x"04", x"04", x"02", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"3C", x"3C", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"3C", x"FF", x"FF", x"FF", x"C3", x"C3", x"E7", x"E7", x"E7", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"02", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"07", x"02", x"02", x"02", x"02", x"02", x"02", x"01", x"00", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"03", x"00", x"00", x"3C", x"C3", x"1C", x"18", x"1C", x"18", x"3C", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"18", x"18", x"3C", x"24", x"18", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"80", x"40", x"40", x"40", x"00", x"00", x"00", x"80", x"C0", x"E0", x"E0", x"E0", x"40", x"40", x"40", x"40", x"40", x"40", x"80", x"00", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"1F", x"3F", x"70", x"60", x"60", x"60", x"60", x"1F", x"20", x"40", x"8F", x"9F", x"98", x"98", x"98", x"60", x"60", x"60", x"60", x"70", x"3F", x"1F", x"00", x"98", x"98", x"98", x"9F", x"8F", x"40", x"20", x"1F", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"F8", x"FC", x"0E", x"06", x"06", x"06", x"06", x"F8", x"04", x"02", x"F1", x"F9", x"19", x"19", x"19", 
															x"06", x"06", x"06", x"06", x"0E", x"FC", x"F8", x"00", x"19", x"19", x"19", x"F9", x"F1", x"02", x"04", x"F8", x"00", x"00", x"00", x"04", x"0A", x"11", x"A0", x"40", x"00", x"00", x"00", x"04", x"0A", x"11", x"A0", x"40", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"38", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"00", x"00", x"00", x"00", x"66", x"7E", x"7E", x"66", x"00", x"00", x"00", x"00", x"00", x"81", x"81", x"00", x"00", x"00", x"00", x"41", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"41", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"40", x"20", x"10", x"08", x"04", x"02", x"01", x"00", x"00", x"00", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"04", x"02", x"01", 
															x"00", x"00", x"00", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"20", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"E0", x"F0", x"38", x"1C", x"0F", x"1F", x"3F", x"3C", x"7F", x"E0", x"00", x"00", x"07", x"1F", x"3C", x"3B", x"00", x"00", x"00", x"00", x"80", x"E0", x"F0", x"F0", x"F8", x"00", x"00", x"00", x"80", x"E0", x"F0", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"1C", x"1C", x"00", x"00", x"07", x"1F", x"3F", x"7C", x"7B", x"7B", x"1F", x"0F", x"58", x"B8", x"33", x"6C", x"E3", x"E0", x"70", x"37", x"E7", x"E7", x"00", x"03", x"E0", x"E0", x"00", x"00", x"00", x"00", x"80", x"E0", x"E0", x"E0", x"00", x"00", x"80", x"E0", x"F0", x"F8", x"78", x"78", 
															x"E0", x"C0", x"60", x"60", x"30", x"D8", x"1C", x"1C", x"38", x"B0", x"80", x"80", x"00", x"00", x"1C", x"1C", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"FF", x"FF", x"81", x"81", x"9D", x"99", x"9D", x"99", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"14", x"14", x"14", x"14", x"14", x"14", x"14", x"14", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"06", x"06", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"39", x"65", x"65", x"65", x"65", x"65", x"39", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"B0", x"B0", x"B6", x"E6", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"04", x"1C", x"B8", x"C0", x"60", x"08", x"14", x"14", x"08", x"00", x"04", x"08", x"F8", x"78", x"7C", x"7C", x"7C", x"3C", x"08", x"00", x"00", x"FE", x"FF", x"7F", x"7F", x"3F", x"1E", x"14", x"08", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E7", x"08", x"14", x"14", x"08", x"08", x"14", x"54", x"2F", x"FF", x"80", x"1F", x"03", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"3F", x"1F", x"0F", x"14", x"08", x"08", x"14", x"84", x"80", x"88", x"F4", x"F4", x"F8", x"08", x"14", x"B4", x"F8", x"C8", x"F4", x"F4", x"F8", x"F8", x"FC", x"FC", x"F8", x"E8", x"D4", x"14", x"08", x"F8", x"FC", x"FC", x"F8", x"E8", x"D4", x"14", x"08", x"10", x"10", x"88", x"80", x"90", x"F0", x"F8", x"F8", x"08", x"08", x"B0", x"FC", x"C8", x"E8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F0", x"F0", x"D0", x"10", x"10", x"F8", x"F8", x"F8", x"F8", x"E8", x"EC", x"6E", x"CA", 
															x"0F", x"1F", x"1E", x"24", x"26", x"70", x"00", x"1F", x"0F", x"1F", x"01", x"1B", x"19", x"0F", x"1F", x"03", x"3F", x"3F", x"7F", x"7E", x"7F", x"3F", x"3C", x"3E", x"00", x"00", x"60", x"7F", x"7F", x"3F", x"04", x"00", x"00", x"E0", x"00", x"80", x"40", x"F0", x"00", x"38", x"00", x"E0", x"80", x"70", x"B8", x"01", x"C3", x"07", x"FC", x"F8", x"E0", x"F4", x"FC", x"F8", x"30", x"00", x"03", x"00", x"20", x"F0", x"F0", x"E0", x"00", x"00", x"00", x"0F", x"1F", x"1E", x"24", x"26", x"70", x"00", x"00", x"0F", x"1F", x"01", x"1B", x"19", x"0F", x"0F", x"1F", x"1F", x"3F", x"7E", x"FF", x"FF", x"C7", x"07", x"18", x"18", x"3C", x"7F", x"7F", x"7F", x"07", x"00", x"00", x"00", x"E0", x"00", x"80", x"40", x"F0", x"00", x"00", x"00", x"E0", x"80", x"70", x"B8", x"00", x"C0", x"80", x"C0", x"E0", x"F0", x"C3", x"C3", x"86", x"C0", x"00", x"00", x"00", x"00", x"BE", x"DE", x"86", x"00", 
															x"1E", x"3F", x"3C", x"49", x"4C", x"E1", x"00", x"39", x"1E", x"3F", x"03", x"36", x"33", x"1E", x"3F", x"3F", x"7F", x"7F", x"7D", x"7F", x"3F", x"1E", x"1C", x"1E", x"00", x"00", x"47", x"7F", x"3F", x"1E", x"00", x"00", x"00", x"C0", x"00", x"00", x"80", x"E0", x"00", x"00", x"08", x"C8", x"04", x"E2", x"71", x"02", x"84", x"08", x"E0", x"E0", x"C0", x"E0", x"E0", x"E0", x"F0", x"00", x"1C", x"1C", x"C8", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"07", x"FF", x"FF", x"3C", x"7F", x"00", x"00", x"00", x"07", x"1F", x"3C", x"3B", x"00", x"00", x"00", x"00", x"80", x"E0", x"F0", x"F0", x"F8", x"00", x"00", x"00", x"80", x"E0", x"F0", x"70", x"00", x"3F", x"7F", x"E0", x"C0", x"C0", x"C1", x"C0", x"C0", x"3F", x"60", x"C0", x"80", x"83", x"8F", x"8F", x"8F", x"D8", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"C7", x"9F", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"87", 
															x"C0", x"C0", x"C0", x"C0", x"C1", x"C3", x"C7", x"C3", x"80", x"80", x"80", x"81", x"83", x"87", x"8F", x"87", x"C1", x"C0", x"C0", x"C0", x"C0", x"E0", x"7F", x"3F", x"81", x"83", x"87", x"8F", x"80", x"C0", x"60", x"3F", x"FF", x"FF", x"01", x"01", x"21", x"11", x"B9", x"43", x"FF", x"00", x"00", x"F0", x"F8", x"FC", x"F8", x"FA", x"03", x"C7", x"97", x"BF", x"7F", x"FF", x"FF", x"FF", x"F2", x"EE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"7D", x"3F", x"7F", x"FD", x"FF", x"FF", x"FF", x"FE", x"7E", x"7E", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"99", x"23", x"01", x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"80", x"80", x"84", x"88", x"9D", x"C2", x"FF", x"00", x"00", x"0F", x"1F", x"3F", x"1F", x"5F", x"C1", x"E1", x"E9", x"FD", x"FE", x"FF", x"FF", x"FF", x"4F", x"77", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", 
															x"FF", x"BE", x"FC", x"FE", x"BF", x"FF", x"FF", x"FF", x"7F", x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"99", x"C4", x"80", x"80", x"80", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"FF", x"FC", x"FE", x"07", x"03", x"03", x"83", x"03", x"03", x"FC", x"06", x"03", x"01", x"C1", x"F1", x"F1", x"F1", x"1B", x"FF", x"FF", x"FF", x"7F", x"FF", x"FF", x"E3", x"F9", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"E1", x"83", x"03", x"03", x"03", x"83", x"C3", x"E3", x"C3", x"81", x"01", x"01", x"81", x"C1", x"E1", x"F1", x"E1", x"83", x"03", x"03", x"03", x"03", x"07", x"FE", x"FC", x"81", x"C1", x"E1", x"F1", x"01", x"03", x"06", x"FC", x"3F", x"7F", x"E0", x"C0", x"C0", x"C0", x"C0", x"C0", x"3F", x"60", x"C0", x"80", x"80", x"80", x"80", x"80", x"C0", x"C7", x"CE", x"DD", x"DF", x"DF", x"DF", x"C7", x"80", x"87", x"8F", x"9F", x"9F", x"9F", x"9F", x"87", 
															x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"0F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"FF", x"FF", x"21", x"C2", x"C0", x"C1", x"E0", x"F1", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"83", x"80", x"9F", x"E0", x"80", x"80", x"E0", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"81", x"01", x"F1", x"0D", x"03", x"02", x"0E", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"F0", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"FF", x"FF", x"8C", x"43", x"03", x"83", x"07", x"8F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"7F", x"FC", x"FE", x"07", x"03", x"03", x"03", x"03", x"03", x"FC", x"06", x"03", x"01", x"01", x"01", x"01", x"01", x"03", x"C3", x"E3", x"33", x"FB", x"FB", x"FB", x"F3", x"01", x"C1", x"E1", x"F1", x"F9", x"F9", x"F9", x"F1", 
															x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"66", x"66", x"66", x"66", x"66", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"19", x"00", x"00", x"03", x"06", x"0C", x"0C", x"18", x"20", x"FF", x"FF", x"00", x"80", x"80", x"80", x"80", x"98", x"00", x"00", x"C0", x"60", x"30", x"30", x"18", x"04", x"00", x"00", x"00", x"00", x"00", x"6C", x"6C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"18", x"04", x"04", x"82", x"42", x"42", x"7E", x"E0", x"F8", x"FC", x"FC", x"FE", x"7E", x"7E", x"7E", x"7F", x"40", x"40", x"40", x"41", x"42", x"42", x"42", x"7F", x"7F", x"7F", x"7F", x"7F", x"7E", x"7E", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"42", x"42", x"42", x"41", x"40", x"40", x"40", x"7F", x"7E", x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"7F", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", 
															x"42", x"43", x"40", x"40", x"40", x"43", x"42", x"42", x"7E", x"7F", x"7F", x"7F", x"7F", x"7F", x"7E", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"42", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"E0", x"18", x"04", x"04", x"82", x"42", x"42", x"42", x"E0", x"F8", x"FC", x"FC", x"FE", x"7E", x"7E", x"7E", x"42", x"42", x"42", x"82", x"04", x"04", x"18", x"E0", x"7E", x"7E", x"7E", x"FE", x"FC", x"FC", x"F8", x"E0", x"7E", x"42", x"42", x"42", x"42", x"42", x"42", x"84", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"FC", x"84", x"08", x"10", x"20", x"10", x"08", x"84", x"84", x"FC", x"F8", x"F0", x"E0", x"F0", x"F8", x"FC", x"FC", x"07", x"18", x"20", x"20", x"41", x"42", x"42", x"42", x"07", x"1F", x"3F", x"3F", x"7F", x"7E", x"7E", x"7E", x"42", x"42", x"42", x"41", x"20", x"20", x"18", x"07", x"7E", x"7E", x"7E", x"7F", x"3F", x"3F", x"1F", x"07", 
															x"FE", x"02", x"02", x"02", x"FE", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"FC", x"04", x"04", x"04", x"FC", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"FE", x"02", x"02", x"02", x"FE", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"78", x"44", x"44", x"42", x"42", x"41", x"41", x"41", x"78", x"7C", x"7C", x"7E", x"7E", x"7F", x"7F", x"7F", x"40", x"40", x"40", x"40", x"40", x"42", x"43", x"43", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"42", x"42", x"42", x"43", x"20", x"20", x"18", x"04", x"7E", x"7E", x"7E", x"7F", x"3F", x"3F", x"1F", x"07", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"C2", x"C2", x"42", x"02", x"02", x"02", x"02", x"02", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", 
															x"82", x"82", x"82", x"42", x"42", x"22", x"22", x"1E", x"FE", x"FE", x"FE", x"7E", x"7E", x"3E", x"3E", x"1E", x"42", x"42", x"42", x"C2", x"04", x"04", x"18", x"20", x"7E", x"7E", x"7E", x"FE", x"FC", x"FC", x"F8", x"E0", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"FF", x"81", x"81", x"81", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"C3", x"42", x"42", x"82", x"02", x"02", x"12", x"EE", x"FF", x"7E", x"7E", x"FE", x"FE", x"FE", x"FE", x"EE", x"00", x"00", x"03", x"0F", x"1F", x"1F", x"3F", x"3F", x"07", x"1F", x"3C", x"70", x"60", x"E0", x"C0", x"C0", x"3F", x"3F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"C0", x"C0", x"E0", x"60", x"70", x"3C", x"1F", x"07", x"00", x"00", x"1F", x"3F", x"3F", x"1F", x"00", x"00", x"3F", x"7F", x"E0", x"C0", x"C0", x"E0", x"7F", x"3F", 
															x"00", x"00", x"80", x"E0", x"E0", x"F0", x"F0", x"F0", x"C0", x"F0", x"78", x"18", x"1C", x"0C", x"0C", x"0C", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F8", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0F", x"07", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"C0", x"C0", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FF", x"FF", x"00", x"00", x"00", x"00", x"03", x"03", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"FC", x"FC", x"F8", x"F8", x"F0", x"C0", x"00", x"00", x"03", x"03", x"07", x"06", x"0E", x"3C", x"F8", x"E0", 
															x"00", x"00", x"F8", x"FC", x"FC", x"F8", x"00", x"00", x"FC", x"FE", x"07", x"03", x"03", x"07", x"FE", x"FC", x"FF", x"FF", x"FE", x"FE", x"FC", x"80", x"80", x"C0", x"00", x"00", x"01", x"01", x"03", x"7F", x"7E", x"30", x"E0", x"E0", x"F0", x"F0", x"E0", x"E0", x"E1", x"E7", x"18", x"1C", x"0C", x"08", x"1B", x"1F", x"1E", x"18", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"3F", x"1F", x"00", x"00", x"01", x"00", x"80", x"C0", x"C0", x"60", x"7F", x"3F", x"06", x"03", x"03", x"07", x"07", x"03", x"83", x"C3", x"F3", x"0C", x"1C", x"18", x"88", x"EC", x"7C", x"3C", x"0C", x"FF", x"7F", x"7F", x"3F", x"3F", x"1F", x"1F", x"0F", x"00", x"80", x"80", x"C0", x"C0", x"E0", x"60", x"70", x"0F", x"07", x"07", x"03", x"03", x"01", x"00", x"00", x"30", x"38", x"18", x"1C", x"0C", x"0E", x"07", x"03", 
															x"00", x"00", x"C0", x"F0", x"F8", x"F8", x"FC", x"FC", x"E0", x"F8", x"3C", x"0E", x"06", x"07", x"03", x"03", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"E0", x"C0", x"C0", x"E0", x"60", x"70", x"30", x"38", x"18", x"E0", x"F0", x"F0", x"E3", x"E7", x"C7", x"CF", x"CF", x"1D", x"0F", x"0F", x"1C", x"18", x"38", x"30", x"30", x"CF", x"CF", x"C7", x"E7", x"E3", x"F0", x"00", x"00", x"30", x"30", x"38", x"18", x"1C", x"0F", x"FF", x"FD", x"0F", x"06", x"06", x"06", x"06", x"06", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"60", x"60", x"66", x"66", x"60", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"99", x"BD", x"A5", x"99", x"81", x"81", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF");
	
	constant SOCCER_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"78", x"FC", x"7C", x"7C", x"FC", x"7C", x"00", x"00", x"78", x"FC", x"0C", x"24", x"04", x"0C", x"60", x"06", x"07", x"01", x"83", x"FF", x"7E", x"7E", x"1C", x"78", x"78", x"7E", x"7C", x"7C", x"7E", x"1E", x"07", x"07", x"06", x"00", x"00", x"00", x"14", x"3C", x"00", x"00", x"08", x"0C", x"0C", x"0C", x"1C", x"3C", x"E2", x"61", x"63", x"21", x"00", x"00", x"00", x"00", x"02", x"1F", x"1F", x"11", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"7C", x"7C", x"FC", x"7C", x"30", x"00", x"78", x"FC", x"0C", x"24", x"04", x"0C", x"0C", x"04", x"0E", x"07", x"1E", x"3E", x"3F", x"3F", x"1E", x"3A", x"30", x"38", x"20", x"26", x"3F", x"27", x"02", x"3B", x"31", x"23", x"01", x"00", x"00", x"14", x"3C", x"07", x"07", x"1B", x"39", x"18", x"18", x"1C", x"3C", x"00", x"D9", x"DD", x"78", x"3E", x"7F", x"FF", x"FF", x"3E", x"26", x"22", x"06", x"0E", x"3F", x"1F", x"08", 
															x"04", x"00", x"00", x"0A", x"1C", x"00", x"00", x"00", x"08", x"0C", x"0C", x"0E", x"1C", x"00", x"00", x"00", x"70", x"30", x"30", x"00", x"00", x"01", x"05", x"0E", x"00", x"00", x"08", x"1C", x"0E", x"07", x"07", x"0E", x"00", x"00", x"78", x"FC", x"FC", x"7C", x"7C", x"7C", x"00", x"00", x"78", x"FC", x"FC", x"04", x"50", x"00", x"00", x"03", x"0B", x"1F", x"3F", x"7F", x"7F", x"F7", x"7F", x"7C", x"74", x"60", x"21", x"3F", x"1C", x"00", x"0E", x"00", x"00", x"00", x"0A", x"1C", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0E", x"1C", x"00", x"00", x"7A", x"32", x"06", x"04", x"00", x"00", x"00", x"00", x"06", x"0E", x"06", x"04", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"FC", x"7C", x"7C", x"7C", x"38", x"00", x"78", x"FC", x"FC", x"04", x"50", x"00", x"06", x"00", x"02", x"03", x"8F", x"FE", x"7E", x"7E", x"7E", x"FE", x"FC", x"FC", x"70", x"70", x"7E", x"30", x"00", 
															x"1E", x"0E", x"0C", x"00", x"01", x"05", x"0E", x"00", x"00", x"00", x"00", x"0E", x"07", x"07", x"0E", x"00", x"03", x"08", x"18", x"18", x"0C", x"03", x"03", x"01", x"00", x"07", x"07", x"07", x"03", x"03", x"03", x"01", x"80", x"08", x"1C", x"0E", x"07", x"F3", x"F2", x"F0", x"70", x"F0", x"E0", x"F0", x"F0", x"F0", x"F0", x"00", x"1E", x"1C", x"00", x"00", x"00", x"30", x"38", x"18", x"00", x"00", x"18", x"18", x"18", x"38", x"38", x"18", x"00", x"78", x"FC", x"FC", x"7C", x"7C", x"78", x"00", x"00", x"78", x"FC", x"FC", x"3C", x"3C", x"18", x"7C", x"20", x"30", x"30", x"18", x"3F", x"7F", x"FF", x"F7", x"5E", x"4E", x"4E", x"66", x"23", x"33", x"1E", x"00", x"FC", x"7E", x"7F", x"7F", x"FF", x"87", x"7E", x"7E", x"1C", x"78", x"78", x"7E", x"78", x"78", x"7E", x"1E", x"30", x"20", x"00", x"02", x"06", x"06", x"04", x"00", x"00", x"18", x"3C", x"1E", x"06", x"06", x"04", x"00", 
															x"00", x"40", x"60", x"60", x"FF", x"FF", x"3F", x"3A", x"7E", x"3E", x"1E", x"1E", x"1F", x"3F", x"1E", x"00", x"3E", x"3E", x"3F", x"3E", x"1C", x"3F", x"3F", x"1E", x"3A", x"30", x"38", x"20", x"22", x"3F", x"27", x"02", x"3E", x"30", x"06", x"06", x"04", x"10", x"38", x"00", x"00", x"04", x"3E", x"1E", x"1C", x"18", x"38", x"00", x"00", x"00", x"78", x"FC", x"FC", x"7C", x"7C", x"78", x"00", x"00", x"78", x"FC", x"FC", x"3C", x"3C", x"18", x"30", x"30", x"2C", x"3C", x"38", x"13", x"03", x"03", x"07", x"0F", x"03", x"03", x"07", x"03", x"03", x"00", x"00", x"18", x"1C", x"0C", x"06", x"F6", x"F4", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"E0", x"38", x"18", x"10", x"00", x"00", x"06", x"06", x"06", x"00", x"00", x"0C", x"0C", x"0E", x"06", x"06", x"06", x"3C", x"7E", x"7E", x"7E", x"7E", x"3C", x"18", x"00", x"3C", x"7E", x"7E", x"42", x"24", x"00", x"67", x"FF", 
															x"40", x"C0", x"C0", x"E0", x"7F", x"3F", x"3F", x"37", x"3F", x"3F", x"3F", x"1F", x"07", x"07", x"3C", x"00", x"3E", x"FF", x"FF", x"7E", x"30", x"7F", x"FF", x"FF", x"3E", x"26", x"22", x"06", x"0E", x"3F", x"1F", x"08", x"66", x"66", x"00", x"00", x"00", x"00", x"05", x"06", x"00", x"10", x"36", x"06", x"06", x"06", x"07", x"06", x"00", x"3C", x"7E", x"7E", x"7E", x"7E", x"3C", x"18", x"00", x"3C", x"7E", x"7E", x"42", x"24", x"00", x"66", x"7F", x"7F", x"7F", x"1F", x"3F", x"7F", x"7F", x"F7", x"7F", x"7C", x"74", x"20", x"21", x"3F", x"1C", x"00", x"00", x"18", x"1C", x"0C", x"38", x"F8", x"E0", x"E0", x"F0", x"E0", x"E0", x"E0", x"C0", x"E0", x"E0", x"80", x"76", x"34", x"00", x"00", x"4A", x"26", x"00", x"00", x"00", x"42", x"66", x"66", x"6E", x"26", x"00", x"00", x"FE", x"FE", x"FF", x"8F", x"FE", x"7E", x"7E", x"7E", x"FE", x"FC", x"FC", x"70", x"70", x"7E", x"30", x"00", 
															x"03", x"0F", x"1F", x"1F", x"0C", x"03", x"03", x"01", x"00", x"07", x"07", x"07", x"03", x"03", x"03", x"01", x"F0", x"F8", x"FC", x"FE", x"07", x"F3", x"F2", x"F0", x"70", x"F0", x"E0", x"F0", x"F0", x"F0", x"F0", x"00", x"7E", x"7E", x"7E", x"18", x"3F", x"7F", x"FF", x"F7", x"5E", x"4E", x"4E", x"66", x"23", x"33", x"1E", x"00", x"1E", x"3F", x"3F", x"3F", x"3F", x"1E", x"00", x"00", x"1E", x"3F", x"3F", x"3F", x"1E", x"0C", x"7E", x"FF", x"30", x"70", x"60", x"37", x"37", x"07", x"06", x"06", x"0F", x"07", x"07", x"07", x"07", x"07", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"E0", x"E0", x"80", x"F0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"60", x"32", x"36", x"06", x"00", x"00", x"00", x"20", x"70", x"07", x"06", x"36", x"30", x"30", x"30", x"30", x"70", x"00", x"3C", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"3C", x"18", x"7E", 
															x"00", x"81", x"81", x"81", x"FF", x"7E", x"7E", x"6E", x"FF", x"7E", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", x"7E", x"7E", x"7E", x"60", x"FF", x"FF", x"3E", x"3A", x"7E", x"3E", x"1E", x"1E", x"1F", x"3F", x"1E", x"00", x"6E", x"00", x"40", x"E4", x"6C", x"0C", x"00", x"00", x"00", x"6C", x"6C", x"EC", x"6C", x"0C", x"00", x"00", x"37", x"3F", x"2F", x"3F", x"38", x"13", x"03", x"03", x"07", x"0F", x"03", x"03", x"03", x"03", x"03", x"00", x"E0", x"F8", x"FC", x"EC", x"06", x"F6", x"F4", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"E0", x"7F", x"FF", x"FF", x"E0", x"7F", x"3F", x"3F", x"37", x"3F", x"3F", x"3F", x"1F", x"07", x"07", x"3C", x"00", x"F0", x"F8", x"FC", x"EC", x"38", x"F8", x"E0", x"E0", x"F0", x"E0", x"E0", x"E0", x"C0", x"E0", x"E0", x"80", x"3F", x"77", x"60", x"37", x"37", x"07", x"06", x"06", x"0F", x"07", x"07", x"07", x"07", x"07", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"78", x"FC", x"7C", x"7C", x"00", x"00", x"00", x"00", x"78", x"FC", x"0C", x"24", x"FC", x"7C", x"10", x"C4", x"FC", x"F8", x"00", x"7C", x"04", x"0C", x"2E", x"3A", x"02", x"06", x"7C", x"7C", x"7C", x"7C", x"F0", x"C0", x"00", x"02", x"56", x"F0", x"7C", x"04", x"00", x"20", x"68", x"6E", x"76", x"F0", x"00", x"00", x"78", x"FC", x"7C", x"7C", x"18", x"E0", x"00", x"00", x"78", x"FC", x"0C", x"24", x"06", x"1F", x"87", x"C0", x"83", x"63", x"01", x"00", x"00", x"00", x"80", x"E0", x"FC", x"7C", x"00", x"00", x"00", x"00", x"F0", x"F0", x"00", x"C2", x"FF", x"79", x"F0", x"E0", x"0C", x"0C", x"FC", x"7C", x"7C", x"38", x"10", x"00", x"18", x"00", x"00", x"00", x"00", x"04", x"0C", x"18", x"00", x"18", x"18", x"1C", x"0C", x"0C", x"0C", x"18", x"F0", x"E0", x"00", x"E0", x"E0", x"E0", x"E0", x"80", x"F0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"60", 
															x"FF", x"FF", x"FF", x"81", x"FF", x"7E", x"7E", x"6E", x"FF", x"7E", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", x"07", x"0F", x"07", x"00", x"00", x"06", x"07", x"07", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"FC", x"03", x"63", x"79", x"1C", x"00", x"00", x"00", x"03", x"00", x"06", x"06", x"03", x"03", x"03", x"03", x"03", x"E0", x"E0", x"84", x"06", x"06", x"0E", x"0C", x"F0", x"20", x"B0", x"78", x"F8", x"F0", x"F0", x"F0", x"F0", x"7E", x"7E", x"78", x"54", x"04", x"08", x"20", x"70", x"7E", x"20", x"00", x"2C", x"3C", x"38", x"30", x"70", x"70", x"78", x"7C", x"FE", x"7C", x"78", x"7C", x"30", x"00", x"00", x"60", x"F0", x"02", x"57", x"07", x"0F", x"80", x"C0", x"C3", x"63", x"03", x"01", x"00", x"00", x"80", x"E0", x"FC", x"7C", x"0C", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"F0", x"F8", x"F8", x"78", x"70", x"FC", x"FC", x"FC", x"FC", x"78", x"78", x"00", x"00", x"C0", x"E0", x"F0", x"F8", x"F8", x"FC", x"E0", x"FC", x"40", x"60", x"F0", x"98", x"98", x"9C", x"1C", x"3C", x"7C", x"FC", x"7E", x"FE", x"FE", x"FE", x"00", x"7C", x"24", x"04", x"0E", x"3A", x"02", x"06", x"7C", x"7C", x"FC", x"FC", x"FC", x"82", x"FF", x"79", x"F0", x"E0", x"0C", x"0C", x"FC", x"7C", x"7C", x"38", x"10", x"00", x"07", x"0F", x"3F", x"7F", x"6F", x"27", x"38", x"1F", x"00", x"0D", x"18", x"0C", x"0F", x"07", x"07", x"07", x"C0", x"E0", x"F8", x"FC", x"EC", x"F8", x"30", x"E0", x"40", x"20", x"70", x"F0", x"E0", x"C0", x"C0", x"E0", x"FC", x"FC", x"0C", x"F0", x"F8", x"F8", x"78", x"70", x"FC", x"FC", x"FC", x"FC", x"78", x"78", x"00", x"00", x"07", x"00", x"00", x"18", x"38", x"70", x"60", x"67", x"03", x"07", x"0F", x"07", x"07", x"07", x"07", x"07", 
															x"C0", x"00", x"00", x"00", x"10", x"10", x"10", x"E0", x"C0", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"7E", x"7E", x"74", x"60", x"00", x"0B", x"1B", x"3A", x"3E", x"1C", x"00", x"12", x"3A", x"1B", x"1B", x"3A", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"7F", x"6C", x"FC", x"C0", x"C4", x"67", x"07", x"03", x"03", x"03", x"83", x"C3", x"FB", x"79", x"09", x"00", x"00", x"00", x"0C", x"0E", x"07", x"F3", x"F3", x"E0", x"80", x"F8", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"00", x"07", x"0F", x"1F", x"1F", x"37", x"38", x"1F", x"07", x"03", x"0F", x"1F", x"07", x"07", x"07", x"07", x"07", x"C0", x"E0", x"F0", x"F8", x"EC", x"1C", x"F8", x"E0", x"C0", x"E0", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"6F", x"FF", x"C3", x"C4", x"67", x"07", x"03", x"03", x"03", x"83", x"C3", x"FB", x"79", x"09", x"00", x"00", 
															x"F8", x"FC", x"FE", x"07", x"F3", x"F3", x"E0", x"80", x"F8", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"00", x"20", x"E0", x"F0", x"F8", x"FC", x"E6", x"0E", x"EC", x"E0", x"40", x"30", x"70", x"E0", x"E0", x"E0", x"E0", x"FC", x"FF", x"E3", x"00", x"E0", x"E0", x"E0", x"E0", x"70", x"F0", x"E0", x"E0", x"E0", x"E0", x"80", x"00", x"E0", x"E0", x"C0", x"80", x"18", x"18", x"0C", x"EC", x"E0", x"C0", x"30", x"70", x"E0", x"E0", x"E0", x"E0", x"FC", x"FC", x"DC", x"88", x"00", x"40", x"D0", x"38", x"FC", x"20", x"00", x"50", x"D8", x"70", x"F0", x"38", x"00", x"00", x"3C", x"7E", x"7E", x"3E", x"7E", x"3C", x"00", x"00", x"3C", x"6E", x"56", x"32", x"34", x"F3", x"24", x"74", x"E4", x"C4", x"C7", x"07", x"07", x"03", x"1F", x"0F", x"07", x"07", x"00", x"00", x"00", x"00", x"8C", x"8F", x"83", x"83", x"E0", x"E0", x"E0", x"E0", x"70", x"F0", x"E0", x"E0", x"E0", x"E0", x"80", x"00", 
															x"E0", x"F0", x"F8", x"FC", x"EC", x"F8", x"18", x"E0", x"E0", x"F0", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"3F", x"FF", x"C7", x"00", x"07", x"07", x"07", x"07", x"0F", x"07", x"07", x"07", x"07", x"07", x"01", x"00", x"FC", x"FF", x"E3", x"00", x"E0", x"C0", x"80", x"00", x"F0", x"E0", x"E0", x"E0", x"E0", x"C0", x"80", x"00", x"FF", x"7E", x"3C", x"42", x"7E", x"7E", x"76", x"76", x"E7", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", x"00", x"66", x"66", x"00", x"00", x"66", x"7E", x"7E", x"00", x"66", x"66", x"66", x"66", x"00", x"3C", x"7E", x"7E", x"62", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"7C", x"FE", x"CC", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"10", x"10", x"18", x"1C", x"EC", x"E0", x"E0", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"FC", x"FC", x"DC", x"CC", x"00", x"00", x"48", x"EC", x"F8", x"70", x"00", x"00", x"CC", x"EC", x"6C", x"EC", 
															x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"30", x"F8", x"C0", x"00", x"07", x"07", x"07", x"07", x"0F", x"07", x"07", x"07", x"07", x"07", x"01", x"00", x"0C", x"1F", x"03", x"00", x"E0", x"C0", x"80", x"00", x"F0", x"E0", x"E0", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"1C", x"1C", x"78", x"FC", x"7C", x"7C", x"00", x"00", x"00", x"00", x"40", x"8C", x"1C", x"4C", x"FC", x"70", x"20", x"00", x"00", x"00", x"00", x"1F", x"44", x"2C", x"1E", x"3E", x"3E", x"3E", x"3F", x"1F", x"00", x"00", x"18", x"3C", x"7C", x"78", x"38", x"38", x"E0", x"F0", x"F8", x"FC", x"FC", x"60", x"00", x"00", x"76", x"76", x"7E", x"7E", x"00", x"7E", x"FF", x"FF", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"FF", x"FF", x"C3", x"81", x"81", x"81", x"BD", x"DB", x"E7", x"66", x"FF", x"7E", x"7E", x"3E", x"00", x"00", x"00", x"00", 
															x"30", x"30", x"30", x"18", x"18", x"0C", x"0F", x"0F", x"00", x"00", x"03", x"07", x"07", x"07", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"FF", x"3A", x"3F", x"3E", x"1C", x"38", x"30", x"30", x"00", x"3D", x"38", x"31", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"07", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"03", x"07", x"04", x"06", x"00", x"00", x"38", x"38", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"C0", x"80", x"90", x"90", x"FF", x"5A", x"00", x"00", x"00", x"00", x"00", x"3F", x"48", x"25", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"78", x"F8", x"F8", x"00", x"00", x"00", x"00", x"00", x"78", x"FE", x"F7", x"7E", x"7E", x"7E", x"00", x"7E", x"7E", x"76", x"76", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"00", x"00", 
															x"76", x"00", x"00", x"00", x"C3", x"C3", x"C3", x"42", x"00", x"66", x"66", x"66", x"E7", x"C3", x"C3", x"42", x"66", x"66", x"E7", x"C3", x"C3", x"81", x"81", x"FF", x"00", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"FF", x"0F", x"1F", x"37", x"7E", x"5C", x"18", x"00", x"00", x"0E", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"80", x"00", x"0E", x"7E", x"7E", x"3E", x"2E", x"38", x"7C", x"FC", x"FE", x"7E", x"7C", x"10", x"00", x"2E", x"00", x"00", x"00", x"00", x"12", x"36", x"6C", x"00", x"36", x"36", x"36", x"36", x"36", x"36", x"6C", x"00", x"00", x"06", x"0F", x"1F", x"3F", x"3F", x"1F", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"03", x"00", x"28", x"74", x"BE", x"54", x"EA", x"54", x"28", x"00", x"38", x"5C", x"EA", x"FE", x"B6", x"7C", x"30", x"00", x"00", x"60", x"F0", x"F0", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"80", x"C0", x"E0", x"E0", x"E0", 
															x"9D", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"FF", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"FF", x"81", x"7E", x"FF", x"FF", x"F7", x"E7", x"24", x"FF", x"FF", x"FF", x"FF", x"99", x"00", x"00", x"C3", x"00", x"00", x"18", x"18", x"18", x"08", x"00", x"00", x"0E", x"0C", x"1C", x"18", x"18", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"33", x"37", x"2F", x"3D", x"1F", x"1F", x"1D", x"08", x"03", x"07", x"0C", x"0A", x"08", x"05", x"02", x"07", x"00", x"00", x"00", x"00", x"00", x"78", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"78", x"FE", x"FF", x"08", x"0C", x"06", x"06", x"0C", x"0C", x"0E", x"0C", x"0F", x"0B", x"01", x"01", x"00", x"00", x"00", x"00", x"EC", x"00", x"00", x"00", x"24", x"6C", x"6C", x"6C", x"00", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", 
															x"C0", x"E0", x"F0", x"B0", x"F8", x"F8", x"B8", x"18", x"C0", x"E0", x"30", x"50", x"18", x"B8", x"48", x"E0", x"00", x"00", x"03", x"00", x"06", x"0F", x"16", x"06", x"07", x"07", x"03", x"0F", x"1F", x"19", x"10", x"00", x"0C", x"0E", x"DD", x"1A", x"09", x"06", x"68", x"60", x"E0", x"E2", x"C3", x"E7", x"FF", x"FE", x"0C", x"00", x"30", x"4B", x"77", x"DF", x"6D", x"3F", x"6F", x"7D", x"28", x"7F", x"BF", x"EC", x"FA", x"58", x"3C", x"1E", x"18", x"08", x"00", x"03", x"00", x"00", x"00", x"06", x"07", x"07", x"07", x"03", x"07", x"0F", x"1F", x"00", x"00", x"00", x"60", x"60", x"F0", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"00", x"C0", x"E0", x"20", x"40", x"BD", x"18", x"00", x"00", x"00", x"00", x"00", x"7E", x"42", x"E7", x"FF", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"F7", x"E7", x"00", x"00", x"42", x"E7", x"7E", x"3C", x"00", x"00", x"C3", x"E7", x"66", x"E7", 
															x"24", x"00", x"81", x"D0", x"C4", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"E0", x"F0", x"F0", x"7E", x"7E", x"BD", x"DB", x"C3", x"C3", x"FF", x"FF", x"FF", x"BD", x"42", x"24", x"3C", x"3C", x"3C", x"18", x"6E", x"66", x"00", x"00", x"00", x"66", x"66", x"42", x"00", x"00", x"66", x"66", x"66", x"66", x"66", x"42", x"33", x"37", x"2F", x"3F", x"1F", x"1F", x"1F", x"08", x"03", x"07", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"C0", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"10", x"C0", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"00", x"00", x"60", x"60", x"F0", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"E0", x"BD", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"FF", x"FF", x"7E", x"7E", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", 
															x"00", x"00", x"81", x"81", x"FF", x"FF", x"FF", x"6E", x"7E", x"FF", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", x"08", x"00", x"03", x"00", x"00", x"00", x"00", x"06", x"07", x"07", x"03", x"07", x"0F", x"1F", x"0F", x"00", x"18", x"1C", x"DE", x"1D", x"0A", x"04", x"18", x"E0", x"E4", x"E2", x"D3", x"E3", x"F7", x"FE", x"FC", x"00", x"10", x"2B", x"57", x"AF", x"5F", x"2F", x"6F", x"77", x"28", x"7F", x"AF", x"FF", x"EF", x"7F", x"3F", x"1F", x"18", x"08", x"00", x"03", x"00", x"00", x"08", x"07", x"07", x"07", x"07", x"03", x"07", x"0F", x"1F", x"07", x"30", x"38", x"78", x"FC", x"7C", x"7C", x"FC", x"64", x"00", x"00", x"60", x"E4", x"24", x"24", x"24", x"3C", x"00", x"40", x"40", x"40", x"FF", x"FF", x"3F", x"33", x"7F", x"3F", x"3F", x"3F", x"3F", x"3F", x"1E", x"00", x"00", x"8C", x"CC", x"DC", x"D8", x"F8", x"F0", x"80", x"00", x"80", x"C0", x"C0", x"40", x"40", x"C0", x"F0", 
															x"C0", x"E0", x"E0", x"FE", x"FE", x"EC", x"C0", x"00", x"C0", x"E0", x"E0", x"80", x"80", x"80", x"78", x"F0", x"03", x"07", x"07", x"03", x"03", x"03", x"01", x"00", x"03", x"07", x"07", x"00", x"02", x"00", x"06", x"0F", x"00", x"00", x"00", x"00", x"00", x"7F", x"FF", x"FF", x"3C", x"3E", x"3E", x"3E", x"3E", x"3F", x"1F", x"08", x"00", x"00", x"00", x"00", x"7C", x"7E", x"3E", x"3C", x"FE", x"7C", x"7C", x"7C", x"7C", x"7E", x"0E", x"04", x"13", x"38", x"78", x"60", x"60", x"03", x"03", x"01", x"0C", x"07", x"07", x"07", x"03", x"03", x"03", x"01", x"60", x"67", x"7F", x"3F", x"1F", x"1F", x"07", x"07", x"00", x"07", x"0F", x"0F", x"00", x"05", x"08", x"0B", x"0C", x"8C", x"DC", x"D8", x"F8", x"F0", x"D0", x"80", x"00", x"80", x"C0", x"C0", x"40", x"00", x"20", x"70", x"30", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"4F", x"7F", x"7F", x"3F", x"3F", x"3F", x"18", x"00", 
															x"88", x"0E", x"0F", x"03", x"03", x"F0", x"F0", x"F0", x"70", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"0C", x"1C", x"78", x"73", x"03", x"03", x"03", x"0F", x"03", x"03", x"03", x"03", x"03", x"01", x"00", x"10", x"18", x"0C", x"0C", x"FC", x"F0", x"E0", x"A0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"E0", x"00", x"30", x"30", x"37", x"1F", x"1F", x"1F", x"17", x"01", x"00", x"00", x"07", x"0F", x"0F", x"03", x"0B", x"0F", x"30", x"30", x"B0", x"E0", x"E0", x"E0", x"E0", x"80", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"E0", x"66", x"66", x"00", x"00", x"00", x"44", x"EE", x"00", x"00", x"00", x"66", x"66", x"66", x"66", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3E", x"FE", x"FE", x"7E", x"7F", x"7F", x"3F", x"3F", x"0E", x"00", x"18", x"1C", x"0E", x"E6", x"E6", x"E0", x"E0", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"80", 
															x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"76", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"1E", x"00", x"C6", x"E6", x"EE", x"EC", x"FC", x"EC", x"C8", x"80", x"C0", x"E0", x"E0", x"20", x"40", x"10", x"B0", x"70", x"20", x"07", x"8F", x"2F", x"07", x"47", x"07", x"03", x"00", x"07", x"0F", x"0F", x"02", x"06", x"02", x"0D", x"00", x"18", x"1C", x"0E", x"E6", x"E6", x"E0", x"60", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"6E", x"68", x"7E", x"7E", x"7E", x"7E", x"7E", x"7C", x"00", x"06", x"C6", x"E6", x"EE", x"EC", x"FC", x"C8", x"00", x"00", x"C0", x"E0", x"E0", x"E0", x"C0", x"B0", x"F0", x"F0", x"04", x"90", x"C5", x"C0", x"F8", x"FA", x"90", x"00", x"00", x"80", x"C0", x"C0", x"00", x"00", x"60", x"F0", x"04", x"00", x"10", x"18", x"0C", x"00", x"00", x"00", x"08", x"0C", x"1C", x"1C", x"0C", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"7C", x"7C", x"FC", x"00", x"00", x"78", x"7C", x"FC", x"0C", x"24", x"04", x"00", x"00", x"00", x"00", x"7C", x"7C", x"FC", x"7C", x"00", x"78", x"7C", x"FC", x"0C", x"24", x"04", x"0C", x"00", x"00", x"00", x"00", x"7C", x"7C", x"7C", x"3E", x"00", x"78", x"7C", x"FC", x"04", x"50", x"00", x"06", x"00", x"00", x"00", x"00", x"00", x"7C", x"7C", x"7C", x"00", x"00", x"78", x"7C", x"FC", x"04", x"50", x"00", x"00", x"00", x"00", x"00", x"7C", x"7C", x"78", x"7C", x"00", x"78", x"7C", x"FC", x"3C", x"3C", x"18", x"7C", x"00", x"00", x"00", x"00", x"00", x"7C", x"7C", x"78", x"00", x"00", x"78", x"7C", x"FC", x"3C", x"3C", x"18", x"00", x"00", x"00", x"42", x"7E", x"3C", x"7F", x"FF", x"3C", x"7E", x"7E", x"7E", x"24", x"00", x"67", x"FF", x"00", x"00", x"00", x"00", x"42", x"7E", x"3C", x"7E", x"00", x"3C", x"7E", x"7E", x"7E", x"24", x"00", x"66", 
															x"00", x"00", x"00", x"3F", x"3F", x"1E", x"7E", x"FF", x"1E", x"3F", x"3F", x"3F", x"1E", x"0C", x"7E", x"FF", x"00", x"00", x"00", x"00", x"7E", x"7E", x"3C", x"7E", x"00", x"3C", x"7E", x"7E", x"7E", x"3C", x"18", x"7E", x"38", x"7C", x"FC", x"FC", x"FE", x"F2", x"30", x"10", x"00", x"0C", x"2A", x"62", x"06", x"0E", x"7C", x"38", x"38", x"7C", x"FE", x"FC", x"F8", x"F6", x"04", x"00", x"20", x"30", x"02", x"1A", x"56", x"CE", x"7C", x"38", x"00", x"00", x"00", x"38", x"7C", x"7C", x"38", x"00", x"00", x"00", x"00", x"38", x"7C", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"00", x"00", x"00", x"00", x"78", x"7C", x"FC", x"0C", x"00", x"00", x"00", x"00", x"7C", x"7C", x"1E", x"FF", x"00", x"78", x"7C", x"FC", x"0C", x"24", x"06", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"FC", 
															x"70", x"78", x"1C", x"0E", x"7E", x"7F", x"7F", x"3F", x"00", x"00", x"60", x"F0", x"02", x"57", x"07", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"7F", x"00", x"00", x"00", x"00", x"10", x"32", x"7E", x"FF", x"00", x"00", x"3C", x"7E", x"7E", x"3E", x"74", x"F3", x"1C", x"3C", x"74", x"E0", x"C7", x"C7", x"07", x"03", x"1F", x"0F", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"1F", x"3F", x"78", x"60", x"00", x"60", x"14", x"38", x"03", x"01", x"00", x"10", x"38", x"78", x"1C", x"38", x"7E", x"7E", x"EE", x"C6", x"00", x"00", x"42", x"E7", x"7C", x"10", x"00", x"00", x"C6", x"67", x"63", x"E7", x"7E", x"F6", x"EE", x"04", x"00", x"00", x"42", x"E7", x"1C", x"00", x"00", x"C2", x"E7", x"63", x"63", x"E7", 
															x"7E", x"7E", x"F7", x"E7", x"81", x"00", x"24", x"E7", x"7E", x"3C", x"00", x"00", x"42", x"E7", x"66", x"E7", x"00", x"66", x"E7", x"C3", x"81", x"81", x"C3", x"FF", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"3C", x"C3", x"34", x"00", x"00", x"10", x"34", x"34", x"00", x"00", x"42", x"76", x"34", x"34", x"34", x"34", x"00", x"00", x"1F", x"1F", x"3F", x"1F", x"0C", x"00", x"00", x"C3", x"03", x"09", x"01", x"03", x"32", x"7F", x"FF", x"FC", x"C7", x"F1", x"F3", x"E3", x"D0", x"C8", x"9C", x"0C", x"F8", x"F0", x"F0", x"60", x"10", x"38", x"7C", x"0C", x"03", x"03", x"07", x"0F", x"8F", x"C1", x"80", x"60", x"03", x"03", x"01", x"00", x"90", x"F8", x"F0", x"60", x"07", x"0F", x"0C", x"08", x"18", x"18", x"3B", x"31", x"07", x"0F", x"0F", x"07", x"07", x"07", x"00", x"00", x"07", x"0F", x"0C", x"08", x"18", x"18", x"3B", x"31", x"07", x"0F", x"0F", x"07", x"07", x"07", x"00", x"00", 
															x"00", x"00", x"1C", x"38", x"30", x"00", x"00", x"02", x"00", x"00", x"1C", x"38", x"38", x"1C", x"0E", x"0C", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"3E", x"3E", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"06", x"2A", x"1E", x"3E", x"30", x"00", x"07", x"0F", x"0F", x"0F", x"01", x"01", x"03", x"03", x"07", x"0F", x"0F", x"01", x"F0", x"60", x"02", x"07", x"03", x"86", x"CE", x"CC", x"08", x"9C", x"FC", x"F8", x"F0", x"E0", x"C0", x"C0", x"1F", x"1F", x"0D", x"83", x"C0", x"C0", x"60", x"00", x"00", x"01", x"31", x"BB", x"F0", x"E0", x"60", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"EC", x"EC", x"F8", x"F8", x"FC", x"FC", x"FC", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"1E", x"3F", x"3F", x"3F", x"3F", x"0E", x"00", x"10", x"1E", x"3F", x"3F", x"1F", x"1F", x"7E", x"FE", x"EE", 
															x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B8", x"9C", x"EE", x"F6", x"F6", x"E0", x"E0", x"80", x"C4", x"E0", x"F0", x"F0", x"F0", x"00", x"00", x"70", x"18", x"1C", x"0C", x"00", x"00", x"00", x"00", x"00", x"78", x"1C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"0F", x"3F", x"70", x"70", x"10", x"00", x"07", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"80", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"E0", x"F0", x"F0", x"00", x"1F", x"1F", x"17", x"07", x"0F", x"07", x"07", x"00", x"07", x"0F", x"00", x"02", x"00", x"06", x"00", x"66", x"00", x"00", x"00", x"88", x"EE", x"66", x"00", x"00", x"66", x"66", x"66", x"EE", x"EE", x"66", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"7E", x"7E", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"42", x"A5", 
															x"11", x"70", x"E0", x"C0", x"07", x"07", x"07", x"07", x"0E", x"0F", x"07", x"07", x"07", x"07", x"07", x"01", x"8E", x"0F", x"03", x"00", x"E0", x"E0", x"E0", x"E0", x"70", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"7A", x"3A", x"38", x"00", x"00", x"30", x"38", x"18", x"00", x"00", x"06", x"38", x"18", x"38", x"38", x"18", x"24", x"00", x"97", x"0F", x"0F", x"30", x"70", x"70", x"00", x"00", x"07", x"0F", x"0F", x"0F", x"0F", x"0F", x"78", x"FC", x"FE", x"5E", x"FF", x"7F", x"23", x"0C", x"78", x"FC", x"8E", x"26", x"07", x"0F", x"1F", x"32", x"00", x"00", x"03", x"00", x"08", x"0C", x"0E", x"0C", x"07", x"07", x"03", x"0F", x"0F", x"03", x"00", x"00", x"E8", x"54", x"BC", x"D2", x"EC", x"74", x"D0", x"E0", x"38", x"FC", x"D6", x"6E", x"BA", x"EC", x"38", x"00", x"07", x"07", x"C7", x"E3", x"E0", x"30", x"18", x"07", x"07", x"07", x"07", x"0F", x"1F", x"0F", x"07", x"07", 
															x"E0", x"E0", x"E0", x"C0", x"0C", x"0E", x"07", x"E3", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"E0", x"E0", x"7C", x"78", x"70", x"3C", x"00", x"10", x"30", x"30", x"7C", x"3C", x"0C", x"0C", x"30", x"30", x"30", x"30", x"00", x"00", x"03", x"00", x"01", x"00", x"07", x"01", x"07", x"07", x"03", x"03", x"07", x"0F", x"0E", x"00", x"D0", x"B8", x"D4", x"FC", x"54", x"E8", x"D0", x"C0", x"70", x"E8", x"7C", x"A8", x"FC", x"B8", x"70", x"00", x"00", x"01", x"02", x"07", x"03", x"05", x"02", x"03", x"03", x"07", x"07", x"05", x"06", x"07", x"07", x"0D", x"C0", x"40", x"E0", x"50", x"B0", x"F0", x"A0", x"40", x"20", x"E0", x"A0", x"F0", x"E0", x"5C", x"F8", x"F0", x"66", x"C3", x"C3", x"81", x"FF", x"C3", x"3C", x"FF", x"00", x"00", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0A", x"00", x"18", x"18", x"18", x"08", x"0F", x"01", x"04", x"0E", x"1C", x"1C", x"18", x"08", 
															x"00", x"00", x"00", x"66", x"66", x"C3", x"C3", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"81", x"FF", x"C3", x"3C", x"FF", x"FF", x"FF", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"08", x"00", x"40", x"00", x"00", x"00", x"00", x"7C", x"7E", x"7E", x"38", x"7C", x"7C", x"7C", x"7C", x"7C", x"7E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"7E", x"7E", x"7E", x"7E", x"FF", x"7E", x"3C", x"18", x"7E", x"66", x"46", x"66", x"E7", x"42", x"3C", x"18", x"7E", x"7E", x"7E", x"7E", x"FF", x"7E", x"3C", x"18", x"7E", x"42", x"7A", x"42", x"CF", x"42", x"3C", x"18", x"18", x"28", x"4F", x"81", x"81", x"4F", x"28", x"18", x"00", x"10", x"30", x"7E", x"7E", x"30", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"C7", x"B3", x"39", x"39", x"39", x"9B", x"C7", x"FF", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"E7", x"C7", x"E7", x"E7", x"E7", x"E7", x"81", x"FF", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"83", x"39", x"F1", x"C3", x"87", x"1F", x"01", x"FF", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"81", x"F3", x"E7", x"C3", x"F9", x"39", x"83", x"FF", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"E3", x"C3", x"93", x"33", x"01", x"F3", x"F3", x"FF", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"03", x"3F", x"03", x"F9", x"F9", x"39", x"83", x"FF", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"C3", x"9F", x"3F", x"03", x"39", x"39", x"83", x"FF", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"01", x"39", x"F3", x"E7", x"CF", x"CF", x"CF", x"FF", 
															x"78", x"C4", x"E4", x"78", x"86", x"86", x"7C", x"00", x"87", x"3B", x"1B", x"87", x"79", x"79", x"83", x"FF", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"83", x"39", x"39", x"81", x"F9", x"F3", x"87", x"FF", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1E", x"06", x"06", x"06", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"AA", x"91", x"AA", x"C4", x"AA", x"11", x"AA", x"44", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"55", x"89", x"55", x"23", x"55", x"88", x"55", x"22", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"7E", x"3C", x"18", x"18", x"18", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"07", x"0F", x"1F", x"3F", x"3F", x"7F", x"7F", x"00", x"00", x"00", x"03", x"07", x"0F", x"0F", x"1F", x"80", x"E0", x"F0", x"F8", x"FC", x"FC", x"FE", x"FE", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"F0", x"F8", 
															x"7F", x"7F", x"3F", x"3F", x"1F", x"0F", x"07", x"01", x"1F", x"0F", x"0F", x"07", x"03", x"00", x"00", x"00", x"FE", x"FE", x"FC", x"FC", x"F8", x"F0", x"E0", x"80", x"F8", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"78", x"78", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"87", x"87", x"FF", x"FF", x"FF", x"00", x"30", x"30", x"00", x"30", x"30", x"00", x"00", x"FF", x"CF", x"CF", x"FF", x"CF", x"CF", x"FF", x"FF", 
															x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"07", x"07", x"02", x"02", x"02", x"02", x"02", x"02", x"04", x"04", x"07", x"07", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"04", x"04", x"04", x"05", x"09", x"0A", x"0A", x"0A", x"0F", x"0F", x"1F", x"1F", x"1F", x"1E", x"1E", x"1E", x"0C", x"0C", x"14", x"14", x"18", x"18", x"19", x"18", x"3E", x"3C", x"3C", x"3C", x"3C", x"38", x"78", x"78", x"31", x"30", x"31", x"32", x"21", x"20", x"65", x"62", x"78", x"70", x"70", x"70", x"F0", x"E0", x"E0", x"E0", x"45", x"48", x"45", x"42", x"85", x"88", x"95", x"82", 
															x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"03", x"03", x"03", x"07", x"01", x"01", x"02", x"02", x"02", x"02", x"02", x"04", x"07", x"07", x"07", x"0F", x"0E", x"0E", x"0E", x"1E", x"04", x"04", x"04", x"08", x"09", x"08", x"09", x"10", x"1C", x"1C", x"1C", x"3C", x"38", x"38", x"38", x"78", x"11", x"12", x"11", x"22", x"25", x"22", x"25", x"42", x"70", x"70", x"70", x"70", x"FA", x"F5", x"EA", x"E0", x"45", x"4A", x"45", x"4A", x"85", x"8A", x"9F", x"8A", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"C0", x"C0", x"95", x"88", x"15", x"22", x"15", x"08", x"15", x"22", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"15", x"08", x"55", x"22", x"55", x"08", x"55", x"22", x"3F", x"7F", x"FF", x"FF", x"C0", x"C0", x"80", x"80", x"7F", x"C0", x"80", x"1F", x"15", x"08", x"55", x"22", 
															x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"55", x"88", x"55", x"22", x"55", x"88", x"55", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"55", x"88", x"55", x"22", x"55", x"88", x"55", x"22", x"00", x"00", x"00", x"00", x"00", x"3F", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"3F", x"40", x"80", x"FF", x"C0", x"C0", x"80", x"80", x"80", x"80", x"80", x"1F", x"28", x"15", x"22", x"55", x"2A", x"55", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"55", x"AA", x"55", x"22", x"55", x"AA", x"55", x"22", x"00", x"00", x"00", x"00", x"AB", x"55", x"AB", x"01", x"55", x"AA", x"55", x"22", x"55", x"AB", x"FF", x"23", x"01", x"01", x"01", x"01", x"01", x"03", x"03", x"03", x"55", x"89", x"55", x"23", x"55", x"8A", x"56", x"22", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"07", x"56", x"8A", x"56", x"22", x"56", x"8A", x"56", x"24", 
															x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"03", x"01", x"FC", x"04", x"04", x"FE", x"56", x"8A", x"56", x"23", x"00", x"00", x"00", x"00", x"00", x"FC", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"FC", x"12", x"12", x"FE", x"1E", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"F2", x"B2", x"61", x"A1", x"61", x"A1", x"65", x"24", x"3F", x"3F", x"3F", x"7F", x"7F", x"7B", x"7B", x"7B", x"64", x"A4", x"64", x"44", x"4C", x"CA", x"4E", x"4A", x"7B", x"7A", x"79", x"79", x"F9", x"F1", x"F1", x"F0", x"4E", x"CA", x"4D", x"4B", x"8D", x"99", x"95", x"92", x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"FF", x"E0", x"95", x"98", x"95", x"92", x"10", x"10", x"3F", x"20", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"C0", x"20", x"20", x"20", x"20", x"20", x"20", x"40", x"40", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", 
															x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"E0", x"E0", x"80", x"80", x"40", x"40", x"40", x"40", x"20", x"20", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"F0", x"20", x"20", x"20", x"10", x"90", x"90", x"90", x"90", x"F9", x"79", x"79", x"79", x"79", x"7D", x"3D", x"3D", x"88", x"C8", x"48", x"48", x"48", x"C4", x"64", x"24", x"3D", x"3D", x"3F", x"1F", x"1F", x"1F", x"1F", x"1F", x"64", x"A4", x"62", x"32", x"52", x"92", x"52", x"31", x"FF", x"FF", x"FF", x"03", x"03", x"03", x"07", x"07", x"09", x"09", x"FF", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"07", x"07", x"06", x"06", x"06", x"86", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"86", x"8E", x"8C", x"8C", x"CC", x"CC", x"CC", x"CC", x"80", x"80", x"80", x"80", x"40", x"40", x"40", x"40", x"CC", x"EC", x"EC", x"EC", x"FC", x"F8", x"F8", x"78", x"40", x"20", x"20", x"20", x"20", x"20", x"10", x"10", 
															x"FF", x"FF", x"F8", x"F8", x"F8", x"F8", x"F8", x"38", x"90", x"90", x"90", x"88", x"48", x"48", x"F8", x"00", x"06", x"06", x"0E", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"0F", x"3F", x"FF", x"3F", x"0F", x"03", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"03", x"03", x"03", x"07", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"70", x"60", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"E0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"06", x"0E", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0C", x"1C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"1F", x"1F", x"18", x"18", x"18", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"F0", x"FC", x"DE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C7", x"C3", x"C1", x"C1", x"C0", x"C0", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"C0", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"81", x"81", x"83", x"83", x"87", x"8E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"BC", x"F8", x"E0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F8", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"38", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"03", x"07", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0C", x"0C", x"0E", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"07", x"03", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0E", x"1C", x"38", x"70", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"70", x"38", x"1C", x"0E", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"1F", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"1F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"3F", x"FF", x"E1", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"07", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"E1", x"FF", x"3F", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"E0", x"40", x"40", x"40", x"40", x"40", x"40", x"20", x"20", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"20", x"20", x"20", x"A0", x"90", x"50", x"50", x"50", x"F0", x"F0", x"F8", x"F8", x"F8", x"78", x"78", x"78", x"30", x"30", x"28", x"28", x"18", x"18", x"98", x"18", 
															x"7C", x"3C", x"3C", x"3C", x"3C", x"1C", x"1E", x"1E", x"8C", x"0C", x"8C", x"4C", x"84", x"04", x"A6", x"46", x"1E", x"0E", x"0E", x"0E", x"0F", x"07", x"07", x"07", x"A2", x"12", x"A2", x"42", x"A1", x"11", x"A9", x"41", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"80", x"80", x"40", x"40", x"40", x"40", x"40", x"20", x"E0", x"E0", x"E0", x"F0", x"70", x"70", x"70", x"78", x"20", x"20", x"20", x"10", x"90", x"10", x"90", x"08", x"38", x"38", x"38", x"3C", x"1C", x"1C", x"1C", x"1E", x"88", x"48", x"88", x"44", x"A4", x"44", x"A4", x"42", x"0E", x"0E", x"0E", x"0E", x"5F", x"AF", x"57", x"07", x"A2", x"52", x"A2", x"52", x"A1", x"51", x"F9", x"51", x"07", x"07", x"07", x"03", x"03", x"03", x"03", x"03", x"A9", x"11", x"A8", x"44", x"A8", x"10", x"A8", x"44", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"A8", x"10", x"AA", x"44", x"AA", x"10", x"AA", x"44", 
															x"FC", x"FE", x"FF", x"FF", x"03", x"03", x"01", x"01", x"FE", x"03", x"01", x"F8", x"A8", x"10", x"AA", x"44", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"11", x"AA", x"44", x"AA", x"11", x"AA", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"11", x"AA", x"44", x"AA", x"11", x"AA", x"44", x"00", x"00", x"00", x"00", x"00", x"FC", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"FC", x"02", x"01", x"FF", x"03", x"03", x"01", x"01", x"01", x"01", x"01", x"F8", x"14", x"A8", x"44", x"AA", x"54", x"AA", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AA", x"55", x"AA", x"44", x"AA", x"55", x"AA", x"44", x"00", x"00", x"00", x"00", x"D5", x"AA", x"D5", x"80", x"AA", x"55", x"AA", x"44", x"AA", x"D5", x"FF", x"C4", x"80", x"80", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"AA", x"91", x"AA", x"C4", x"AA", x"51", x"6A", x"44", 
															x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"6A", x"51", x"6A", x"44", x"6A", x"51", x"6A", x"24", x"FF", x"FF", x"FF", x"FF", x"C0", x"C0", x"C0", x"80", x"3F", x"20", x"20", x"7F", x"6A", x"51", x"6A", x"C4", x"00", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"3F", x"48", x"48", x"7F", x"78", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"4F", x"4D", x"86", x"85", x"86", x"85", x"A6", x"24", x"FC", x"FC", x"FC", x"FE", x"FE", x"DE", x"DE", x"DE", x"26", x"25", x"26", x"22", x"32", x"53", x"72", x"52", x"DE", x"5E", x"9E", x"9E", x"9F", x"8F", x"8F", x"0F", x"72", x"53", x"B2", x"D2", x"B1", x"99", x"A9", x"49", x"0F", x"0F", x"0F", x"0F", x"FF", x"FF", x"FF", x"07", x"A9", x"19", x"A9", x"49", x"08", x"08", x"FC", x"04", x"07", x"07", x"07", x"07", x"07", x"07", x"03", x"03", x"04", x"04", x"04", x"04", x"04", x"04", x"02", x"02", 
															x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"03", x"03", x"03", x"03", x"07", x"07", x"01", x"01", x"02", x"02", x"02", x"02", x"04", x"04", x"07", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"0F", x"04", x"04", x"04", x"08", x"09", x"09", x"09", x"09", x"9F", x"9E", x"9E", x"9E", x"9E", x"BE", x"BC", x"BC", x"11", x"13", x"12", x"12", x"12", x"23", x"26", x"24", x"BC", x"BC", x"FC", x"F8", x"F8", x"F8", x"F8", x"F8", x"26", x"25", x"46", x"4C", x"4A", x"49", x"4A", x"8C", x"FF", x"FF", x"FF", x"C0", x"C0", x"C0", x"E0", x"E0", x"90", x"90", x"FF", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"E0", x"E0", x"60", x"60", x"60", x"61", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"61", x"71", x"31", x"31", x"33", x"33", x"33", x"33", x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"02", 
															x"33", x"37", x"37", x"37", x"3F", x"1F", x"1F", x"1E", x"02", x"04", x"04", x"04", x"04", x"04", x"08", x"08", x"FF", x"FF", x"1F", x"1F", x"1F", x"1F", x"1F", x"1C", x"09", x"09", x"09", x"11", x"12", x"12", x"1F", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"F0", x"FC", x"FF", x"FC", x"F0", x"C0", x"C0", x"C0", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0E", x"06", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"06", x"06", x"06", x"07", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"60", x"70", x"30", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"30", x"38", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"F8", x"F8", x"18", x"18", x"18", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"06", x"06", x"06", x"0F", x"3F", x"7B", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E3", x"C3", x"83", x"83", x"03", x"03", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"03", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"81", x"81", x"C1", x"C1", x"E1", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3D", x"1F", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"1C", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"06", x"06", x"06", x"06", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"03", x"03", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"C0", x"E0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"70", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"30", x"30", x"70", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"E0", x"C0", x"C0", x"C0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"70", x"38", x"1C", x"0E", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"07", x"0E", x"1C", x"38", x"70", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F8", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"F8", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"FC", x"FF", x"87", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"80", x"87", x"FF", x"FC", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"06", x"0E", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"1C", x"18", x"18", x"1C", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1B", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"38", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"30", x"30", x"30", x"70", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"60", x"60", x"60", x"E0", x"C0", x"C0", x"C3", x"CF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"F8", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"60", x"60", x"60", x"70", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"38", x"18", x"18", x"18", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"D8", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"1C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0E", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"06", x"06", x"06", x"07", x"03", x"03", x"C3", x"F3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"1F", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"03", x"03", x"03", x"03", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"00");
	
	constant F1_RACE_CHR_ROM : CHR_ROM_ARRAY := (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"1F",x"16",x"00",x"00",x"0C",x"0B",x"0B",x"0C",x"0C",x"03",x"77",x"E7",x"CE",x"FF",x"FF",x"FF",x"FF",x"07",x"7E",x"FC",x"31",x"FF",x"FF",x"00",x"03",
																x"00",x"00",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"5E",x"00",x"00",x"00",x"E1",x"E3",x"E7",x"C7",x"8F",x"BF",x"FF",x"BF",x"DE",x"DD",x"DB",x"BB",x"70",x"49",x"05",x"4C",x"FF",x"3C",x"BD",x"BD",x"FF",x"FF",x"FF",x"FF",x"3C",x"FF",x"FF",x"7E",x"3C",x"5A",x"66",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"FF",x"FC",x"BC",x"E7",x"B5",x"9F",x"80",x"00",x"00",x"03",x"13",x"00",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"00",x"24",x"24",x"18",x"E7",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"10",x"10",x"10",x"10",x"10",x"38",x"38",x"38",x"00",x"00",x"00",x"00",x"00",
																x"00",x"08",x"3C",x"28",x"00",x"10",x"10",x"10",x"7C",x"7C",x"7C",x"7C",x"7C",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"1F",x"1F",x"1F",x"9F",x"FF",x"FF",x"FF",x"F1",x"0B",x"00",x"00",x"80",x"7F",x"7F",x"80",x"EE",
																x"83",x"87",x"B7",x"CC",x"FF",x"FF",x"FF",x"FF",x"03",x"06",x"0C",x"33",x"FF",x"FF",x"00",x"70",x"E0",x"F1",x"F1",x"6D",x"FC",x"FC",x"FC",x"0C",x"DC",x"6F",x"2F",x"96",x"F7",x"F7",x"07",x"F7",x"3F",x"BF",x"FF",x"FF",x"BF",x"3F",x"3F",x"9E",x"1A",x"80",x"C0",x"00",x"00",x"00",x"80",x"C0",x"01",x"01",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"5E",x"00",x"00",x"00",
																x"F3",x"E6",x"E7",x"CF",x"DF",x"FF",x"FF",x"DF",x"EC",x"DB",x"DB",x"B1",x"28",x"02",x"0A",x"39",x"FF",x"79",x"7B",x"7B",x"FF",x"FF",x"FF",x"FF",x"78",x"FF",x"FF",x"FD",x"78",x"B5",x"CD",x"FE",x"8C",x"8C",x"EF",x"FF",x"F7",x"FF",x"FF",x"F7",x"77",x"77",x"B4",x"90",x"2B",x"00",x"40",x"68",x"80",x"00",x"FC",x"FF",x"FF",x"FE",x"FF",x"FE",x"C0",x"C0",x"00",x"00",x"D0",x"04",x"04",x"04",
																x"FF",x"F9",x"F9",x"EF",x"BB",x"9F",x"80",x"00",x"00",x"06",x"26",x"01",x"02",x"00",x"00",x"00",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF",x"FC",x"00",x"48",x"49",x"31",x"CE",x"79",x"78",x"00",x"00",x"FF",x"7F",x"77",x"DF",x"77",x"E7",x"07",x"03",x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",
																x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"00",x"00",x"00",x"F0",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"F0",x"BF",x"BF",x"C0",x"E0",x"3F",x"3F",x"3F",x"3F",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"C0",x"8F",x"9F",x"A1",x"7F",x"FF",x"FF",x"FF",x"BF",x"0F",x"39",x"5E",x"9C",x"DE",x"DE",x"1E",x"5E",x"C0",x"E7",x"E7",x"E3",x"C2",x"C0",x"80",x"04",x"30",x"9F",x"9F",x"1C",x"3C",x"3C",x"7E",x"FE",
																x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"7C",x"70",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"2E",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"EF",x"FF",x"FF",x"BF",x"F9",x"FB",x"F7",x"E3",x"10",x"05",x"15",x"73",x"FF",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E6",x"FE",x"FF",x"FB",x"F0",x"6A",x"9A",x"FC",
																x"3E",x"3C",x"BF",x"BF",x"9F",x"DF",x"FF",x"DF",x"DF",x"DF",x"58",x"40",x"67",x"20",x"80",x"E0",x"08",x"00",x"F8",x"FC",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"06",x"00",x"40",x"08",x"0C",x"0C",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"F3",x"F3",x"FF",x"EF",x"CF",x"01",x"00",x"40",x"2C",x"2C",x"03",x"04",x"00",x"00",x"00",
																x"FF",x"FC",x"FC",x"FF",x"FE",x"FF",x"F8",x"00",x"90",x"93",x"63",x"9C",x"F2",x"F0",x"00",x"00",x"FF",x"FF",x"FF",x"9F",x"FF",x"9F",x"0F",x"07",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FC",x"F8",x"0C",x"0C",x"0C",x"0C",x"04",x"00",x"00",x"00",x"1F",x"3F",x"3E",x"3C",x"00",x"00",x"03",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
																x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"1F",x"00",x"16",x"00",x"0C",x"0B",x"0B",x"0C",x"0C",x"00",x"00",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"5E",x"5E",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"1F",x"1F",x"9F",x"FF",x"FF",x"FF",x"F1",x"00",x"0B",x"00",x"80",x"7F",x"7F",x"80",x"EE",
																x"FC",x"38",x"30",x"20",x"00",x"00",x"C0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"3F",x"BF",x"FF",x"FF",x"BF",x"3F",x"3F",x"9E",x"00",x"9A",x"C0",x"00",x"00",x"00",x"80",x"C0",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"00",x"5E",x"5E",x"00",x"8C",x"8C",x"EF",x"CF",x"D7",x"FF",x"FF",x"F7",x"77",x"77",x"B4",x"B0",x"28",x"03",x"43",x"68",
																x"80",x"00",x"FC",x"FE",x"FE",x"FE",x"FE",x"FE",x"C0",x"C0",x"00",x"00",x"00",x"D4",x"D4",x"04",x"FF",x"1F",x"8F",x"FF",x"1F",x"8F",x"8F",x"1F",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"3F",x"3F",x"3F",x"3F",x"FF",x"FF",x"FF",x"FF",x"1C",x"00",x"00",x"00",x"FF",x"FF",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"7C",x"00",x"74",x"04",x"04",x"04",x"04",x"00",x"00",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"5C",x"5C",x"00",x"00",x"00",x"3E",x"3C",x"FF",x"BF",x"9F",x"DF",x"FF",x"DF",x"DF",x"DF",x"58",x"40",x"60",x"2E",x"8E",x"E0",x"08",x"00",x"F8",x"FC",x"FF",x"FE",x"FF",x"FE",x"FF",x"FE",x"06",x"00",x"00",x"88",x"8C",x"0C",
																x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"DB",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"E7",x"07",x"07",x"07",x"03",x"01",x"7D",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"5C",x"E2",x"FF",x"FF",x"FF",x"C9",x"DD",x"9D",x"3F",x"8D",x"7F",x"7F",x"80",x"B7",x"AF",x"63",x"C5",
																x"FE",x"FE",x"FF",x"FF",x"FF",x"FE",x"FE",x"7C",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"E7",x"E7",x"BF",x"EB",x"7F",x"00",x"16",x"43",x"1A",x"19",x"06",x"03",x"01",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"7C",x"5D",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"03",x"1F",x"3F",x"73",x"62",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"3B",x"65",x"00",x"00",x"00",x"00",x"00",x"0E",x"DF",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"CC",x"E0",x"03",x"03",x"03",x"03",x"03",x"7F",x"FF",x"FF",x"03",x"02",x"02",x"03",x"03",x"03",x"02",x"58",
																x"7C",x"FF",x"FF",x"FF",x"8F",x"93",x"3B",x"3F",x"01",x"FF",x"FF",x"00",x"72",x"6F",x"DF",x"C3",x"4E",x"FE",x"FE",x"FE",x"C6",x"36",x"77",x"FB",x"B3",x"FB",x"FB",x"03",x"3B",x"CB",x"EA",x"04",x"7F",x"1F",x"1F",x"0E",x"00",x"FC",x"FE",x"FE",x"80",x"80",x"C0",x"E0",x"E0",x"00",x"00",x"D0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"FF",x"FF",x"4F",x"CF",x"BF",x"D7",x"7F",x"00",x"2C",x"07",x"B4",x"33",x"0C",x"07",x"03",x"00",x"FF",x"FB",x"CF",x"CF",x"F7",x"AD",x"F9",x"00",x"D0",x"86",x"B0",x"30",x"C0",x"80",x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"7C",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"58",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"D4",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"1E",x"3F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"85",
																x"00",x"00",x"00",x"00",x"00",x"1E",x"3F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"82",x"03",x"03",x"03",x"03",x"7F",x"FF",x"FF",x"FF",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"58",x"C3",x"FF",x"FF",x"FF",x"FF",x"C6",x"B6",x"7F",x"C0",x"7F",x"7F",x"80",x"84",x"BF",x"4F",x"86",x"CF",x"FF",x"FF",x"FF",x"FE",x"4F",x"EF",x"E7",x"37",x"F7",x"F7",x"07",x"07",x"B6",x"D4",x"19",
																x"E7",x"C3",x"8B",x"11",x"00",x"FC",x"FE",x"FE",x"18",x"38",x"7C",x"FC",x"F8",x"00",x"00",x"A0",x"F0",x"F0",x"F0",x"E0",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"9F",x"FF",x"AF",x"7F",x"00",x"59",x"8F",x"69",x"66",x"19",x"0F",x"06",x"00",
																x"DB",x"FB",x"9F",x"9B",x"EF",x"4B",x"FB",x"01",x"A4",x"04",x"68",x"60",x"80",x"00",x"00",x"00",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"04",x"0C",x"0C",x"0C",x"04",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"58",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"DB",x"FB",x"9F",x"9B",x"E7",x"4B",x"FB",x"01",x"A5",x"04",x"68",x"60",x"80",x"00",x"00",x"00",
																x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"A4",x"0C",x"0C",x"0C",x"04",x"00",x"00",x"00",x"00",x"00",x"0E",x"0E",x"0F",x"0F",x"0F",x"06",x"00",x"00",x"00",x"00",x"04",x"07",x"06",x"05",x"00",x"00",x"24",x"DB",x"BD",x"FF",x"FF",x"3C",x"00",x"00",x"3C",x"FF",x"42",x"FF",x"00",x"DB",x"FF",x"F8",x"FF",x"FF",x"FE",x"FB",x"F9",x"F8",x"05",x"B3",x"04",x"00",x"00",x"00",x"00",x"00",
																x"5A",x"DB",x"FF",x"7E",x"FF",x"7E",x"FF",x"00",x"FF",x"3C",x"24",x"99",x"66",x"3C",x"18",x"00",x"00",x"00",x"00",x"00",x"06",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"06",x"05",x"06",x"06",x"00",x"00",x"00",x"E3",x"F1",x"FF",x"FF",x"7C",x"00",x"00",x"00",x"03",x"0E",x"FF",x"00",x"B3",x"00",x"00",x"00",x"0E",x"AE",x"9E",x"8E",x"80",x"00",x"00",x"00",x"C0",x"C0",x"E0",x"E0",x"F0",
																x"7C",x"FC",x"FD",x"FE",x"FD",x"FE",x"FD",x"78",x"0F",x"03",x"E2",x"01",x"00",x"00",x"00",x"00",x"B5",x"B4",x"FF",x"FD",x"FE",x"FD",x"FF",x"00",x"FE",x"7B",x"48",x"32",x"CC",x"78",x"30",x"00",x"BC",x"FF",x"7E",x"FE",x"FE",x"7E",x"7E",x"3C",x"C0",x"00",x"74",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"E3",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"E0",x"BF",x"C0",
																x"00",x"00",x"00",x"C0",x"CE",x"BF",x"FE",x"F8",x"00",x"00",x"00",x"00",x"15",x"5A",x"59",x"1F",x"00",x"00",x"00",x"1E",x"1E",x"3E",x"1E",x"1E",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"E0",x"7F",x"FF",x"FD",x"FB",x"FA",x"FD",x"FF",x"7C",x"0E",x"0C",x"72",x"04",x"05",x"00",x"00",x"00",x"63",x"6B",x"6C",x"FF",x"F6",x"FB",x"FE",x"00",x"FD",x"FD",x"F3",x"90",x"09",x"F0",x"60",x"00",
																x"FC",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"7C",x"80",x"00",x"74",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"1F",x"3F",x"00",x"00",x"00",x"00",x"00",x"1E",x"18",x"1C",x"00",x"00",x"00",x"00",x"00",x"1F",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"0F",x"EF",x"0F",x"00",x"00",x"00",x"00",x"38",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"48",x"F6",x"F3",x"FF",
																x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C4",x"7F",x"7E",x"7C",x"7B",x"7B",x"7F",x"3C",x"00",x"1E",x"2D",x"03",x"06",x"05",x"01",x"00",x"00",x"FF",x"CF",x"C7",x"F7",x"FF",x"FF",x"F7",x"03",x"8C",x"F8",x"FB",x"18",x"20",x"E0",x"C0",x"00",x"F5",x"FA",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"0F",x"07",x"27",x"77",x"74",x"20",x"00",x"00",
																x"3E",x"1E",x"1C",x"00",x"00",x"00",x"00",x"00",x"C4",x"C4",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3A",x"3D",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"12",x"03",x"01",x"1F",x"1E",x"1F",x"1F",x"1E",x"1E",x"01",x"01",x"01",x"17",x"00",x"00",x"00",x"00",x"FF",x"FF",x"99",x"3C",x"FF",x"5A",x"FF",x"00",x"FF",x"18",x"7E",x"C3",x"18",x"24",x"18",x"00",
																x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"37",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"03",x"03",x"1E",x"1E",x"1E",x"1F",x"1E",x"1E",x"03",x"03",x"01",x"1D",x"00",x"00",x"00",x"00",x"FF",x"FF",x"B5",x"CE",x"7A",x"FB",x"FE",x"00",x"FF",x"31",x"CF",x"31",x"CC",x"78",x"30",x"00",
																x"70",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"80",x"C0",x"00",x"E0",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E4",x"EE",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"15",x"00",x"00",x"00",x"00",x"00",x"00",x"70",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"1F",x"0F",x"7C",x"FB",x"FD",x"FF",x"FB",x"70",x"1F",x"0C",x"0B",x"64",x"02",x"01",x"00",x"00",x"F8",x"F8",x"97",x"EF",x"DF",x"FF",x"EF",x"07",x"DF",x"9F",x"F8",x"16",x"A1",x"41",x"80",x"00",x"F0",x"70",x"00",x"80",x"80",x"80",x"80",x"00",x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3A",x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"3F",x"79",x"77",x"7F",x"7F",x"3B",x"00",x"1F",x"19",x"17",x"08",x"02",x"03",x"01",x"00",x"F3",x"F0",x"3E",x"BF",x"FF",x"FF",x"BF",x"1E",x"FD",x"3F",x"E1",x"40",x"82",x"82",x"00",x"00",
																x"0E",x"0E",x"0E",x"0E",x"00",x"00",x"00",x"00",x"C0",x"F2",x"F2",x"E0",x"80",x"00",x"00",x"00",x"00",x"00",x"20",x"30",x"38",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"18",x"1F",x"09",x"73",x"77",x"79",x"77",x"70",x"03",x"0F",x"0F",x"0D",x"08",x"02",x"01",x"00",x"03",x"0F",x"0F",x"7B",x"77",x"7D",x"77",x"70",x"00",x"0C",x"0F",x"0D",x"09",x"02",x"01",x"00",
																x"06",x"16",x"F0",x"9E",x"CE",x"BE",x"EE",x"0E",x"70",x"F8",x"F8",x"70",x"30",x"40",x"80",x"00",x"00",x"0F",x"0F",x"7D",x"73",x"7F",x"77",x"70",x"00",x"0F",x"0D",x"0B",x"04",x"02",x"01",x"00",x"C3",x"F3",x"E3",x"3C",x"9C",x"FC",x"DC",x"1C",x"00",x"EC",x"3C",x"E0",x"60",x"80",x"00",x"00",x"00",x"01",x"01",x"07",x"0F",x"0F",x"0F",x"07",x"00",x"01",x"01",x"01",x"00",x"01",x"00",x"00",
																x"00",x"FD",x"FC",x"AF",x"6F",x"FF",x"6F",x"07",x"00",x"FE",x"AF",x"78",x"91",x"61",x"01",x"00",x"00",x"00",x"8C",x"0C",x"8C",x"80",x"80",x"00",x"00",x"00",x"40",x"F0",x"70",x"40",x"00",x"00",x"00",x"00",x"00",x"04",x"07",x"19",x"1D",x"1A",x"00",x"00",x"00",x"01",x"07",x"07",x"02",x"03",x"00",x"00",x"00",x"03",x"07",x"1B",x"1F",x"1B",x"00",x"00",x"00",x"00",x"07",x"05",x"02",x"01",
																x"00",x"00",x"00",x"18",x"C0",x"98",x"F8",x"D8",x"00",x"00",x"00",x"E0",x"E0",x"60",x"40",x"80",x"00",x"00",x"00",x"03",x"0F",x"32",x"3F",x"37",x"00",x"00",x"00",x"00",x"0F",x"07",x"05",x"06",x"00",x"00",x"00",x"18",x"98",x"60",x"E0",x"60",x"00",x"00",x"00",x"40",x"E0",x"80",x"00",x"00",x"00",x"00",x"00",x"0F",x"04",x"36",x"3F",x"36",x"00",x"00",x"00",x"0F",x"07",x"09",x"04",x"00",
																x"00",x"00",x"00",x"40",x"06",x"E6",x"E0",x"E0",x"00",x"00",x"00",x"C0",x"F0",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"3C",x"3C",x"24",x"00",x"00",x"00",x"00",x"00",x"38",x"52",x"5A",x"00",x"00",x"00",x"00",x"00",x"3E",x"3C",x"24",x"00",x"00",x"00",x"00",x"00",x"39",x"D6",x"D6",x"00",x"00",x"00",x"00",x"00",x"3E",x"38",x"28",
																x"00",x"00",x"00",x"00",x"00",x"71",x"ED",x"CC",x"00",x"00",x"00",x"00",x"00",x"7C",x"32",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"01",x"82",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"01",x"00",x"00",x"00",x"00",x"04",x"01",x"02",
																x"01",x"07",x"1D",x"33",x"7E",x"DD",x"BF",x"FF",x"01",x"37",x"7E",x"BC",x"69",x"E2",x"C0",x"00",x"FF",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"01",x"04",x"00",x"01",x"00",x"EF",x"FF",x"F7",x"F9",x"5F",x"2F",x"1E",x"03",x"10",x"00",x"88",x"C6",x"E0",x"30",x"3D",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"30",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"30",x"70",x"70",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"38",x"1F",x"0F",x"07",x"03",x"E1",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"3D",x"1D",x"1F",x"DF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"20",x"F0",x"F0",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"E0",x"E0",x"C0",x"C0",x"C0",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"0F",x"07",x"03",x"0F",x"3F",x"1F",x"0F",x"00",x"20",x"06",x"0B",x"0F",x"3F",x"3F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"F8",x"00",x"C0",x"E9",x"BC",x"FC",x"F8",x"FE",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"2F",x"9F",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"F8",x"F0",x"E0",x"FC",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"0F",x"1F",x"7F",x"FF",x"03",x"00",x"00",x"7D",x"3F",x"1F",x"3F",x"3F",x"1F",x"0F",x"07",x"F2",x"F0",x"F8",x"F2",x"F0",x"F8",x"F8",x"DC",x"FF",x"DE",x"FA",x"FE",x"FC",x"FC",x"F8",x"F0",x"07",x"27",x"0F",x"07",x"0F",x"2F",x"1F",x"3E",
																x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"F8",x"F0",x"E0",x"F0",x"F8",x"FC",x"9E",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"00",x"60",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"06",x"07",x"03",x"03",x"03",x"21",x"19",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"98",x"9C",x"CE",x"EE",x"F7",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"40",x"40",x"C3",x"C7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"03",x"07",x"1F",x"3E",x"7C",x"FC",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"40",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"30",x"00",x"03",x"01",x"00",x"00",
																x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"1F",x"0F",x"0F",x"07",x"07",x"E7",x"7B",x"7F",x"00",x"00",x"10",x"0C",x"06",x"67",x"35",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"07",x"8F",x"DE",x"BC",x"CF",x"DF",x"EF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"00",x"00",x"00",x"C0",x"C0",x"80",x"F0",x"F8",x"FC",x"F8",x"F0",x"F8",x"FF",x"FF",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"1C",x"F8",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"03",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"01",x"07",x"03",x"03",x"01",x"01",x"03",x"3F",x"FF",x"FF",x"7F",x"3F",x"7F",x"3F",x"0F",x"7F",x"FF",x"E7",x"AF",x"FF",x"FF",x"7F",x"F7",x"FF",x"FC",x"F8",x"F0",x"C1",x"C2",x"E0",x"C8",
																x"FB",x"FD",x"FC",x"FE",x"E7",x"F7",x"FF",x"FF",x"FF",x"E3",x"43",x"21",x"18",x"09",x"00",x"00",x"C0",x"80",x"B8",x"F8",x"F0",x"F0",x"B8",x"DC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"E0",x"C0",x"80",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"00",x"00",x"00",x"00",
																x"07",x"07",x"03",x"01",x"00",x"01",x"00",x"00",x"3F",x"FF",x"FF",x"FF",x"3F",x"03",x"07",x"00",x"FF",x"FF",x"7F",x"B7",x"F3",x"FF",x"FF",x"3F",x"00",x"80",x"A0",x"C8",x"CC",x"80",x"E2",x"3C",x"FF",x"FF",x"FF",x"FF",x"FE",x"F7",x"FF",x"FF",x"02",x"02",x"04",x"00",x"01",x"0A",x"00",x"31",x"FB",x"FF",x"F8",x"70",x"E0",x"E0",x"C0",x"00",x"FF",x"7F",x"3F",x"9F",x"3E",x"7F",x"E7",x"80",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"F8",x"FF",x"C0",x"00",x"00",x"C0",x"00",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"38",x"00",x"00",x"38",x"38",x"38",x"00",x"00",x"00",x"38",x"38",x"38",x"38",x"38",x"38",x"38",
																x"38",x"38",x"38",x"00",x"00",x"00",x"00",x"00",x"38",x"38",x"38",x"38",x"38",x"38",x"00",x"00",x"38",x"7C",x"04",x"08",x"04",x"4C",x"7C",x"7C",x"00",x"00",x"78",x"74",x"78",x"74",x"78",x"74",x"7C",x"7C",x"3C",x"08",x"04",x"08",x"44",x"7C",x"78",x"74",x"78",x"74",x"78",x"74",x"78",x"74",x"7C",x"7C",x"7C",x"38",x"04",x"08",x"04",x"08",x"78",x"74",x"78",x"74",x"78",x"74",x"78",x"30",
																x"7E",x"FF",x"7E",x"05",x"02",x"05",x"02",x"85",x"00",x"00",x"81",x"FA",x"FD",x"FA",x"FD",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FD",x"FA",x"FD",x"FA",x"FD",x"FA",x"FD",x"FA",x"02",x"05",x"02",x"05",x"02",x"05",x"02",x"85",x"FD",x"FA",x"FD",x"FA",x"FD",x"FA",x"FD",x"FA",x"02",x"05",x"02",x"05",x"02",x"05",x"02",x"04",x"FD",x"FA",x"FD",x"FA",x"FD",x"FA",x"FD",x"7A",
																x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"38",x"28",x"38",x"28",x"38",x"38",x"38",x"00",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"00",x"7E",x"66",x"66",x"7E",x"66",x"66",x"7E",x"66",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"7E",x"6E",x"66",x"7E",x"7E",x"7E",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",
																x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"C7",x"9F",x"93",x"C3",x"FF",x"C7",x"93",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"93",x"C7",x"FF",x"C7",x"93",x"83",x"93",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"9F",x"9F",x"9F",x"83",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",
																x"FF",x"F8",x"F0",x"F1",x"F1",x"F1",x"F1",x"F8",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"1F",x"0F",x"8F",x"FF",x"0F",x"8F",x"0F",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FF",x"FC",x"F8",x"F1",x"F1",x"F0",x"F0",x"F1",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"F1",x"F1",x"F1",x"F1",x"F1",x"F0",x"F0",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"0F",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"7E",x"7E",x"7E",x"66",x"66",x"7E",x"66",x"66",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"9F",x"93",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"C3",x"FF",x"C7",x"93",x"93",x"C7",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"F8",x"F1",x"F1",x"F8",x"FF",x"F1",x"F8",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",
																x"FF",x"F0",x"F0",x"FE",x"FE",x"FE",x"FE",x"FE",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"F0",x"F1",x"F1",x"F0",x"F1",x"F1",x"F1",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"1F",x"8F",x"8F",x"1F",x"3F",x"9F",x"CF",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"09",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"09",
																x"00",x"00",x"00",x"00",x"20",x"80",x"D8",x"A4",x"00",x"00",x"00",x"00",x"20",x"80",x"D8",x"A4",x"00",x"02",x"00",x"01",x"0A",x"1F",x"36",x"20",x"00",x"02",x"00",x"01",x"0A",x"1F",x"36",x"20",x"00",x"00",x"00",x"C0",x"E0",x"D8",x"BC",x"22",x"00",x"00",x"00",x"C0",x"E0",x"D8",x"BC",x"22",x"06",x"1F",x"3B",x"75",x"5A",x"15",x"00",x"00",x"06",x"1F",x"3B",x"75",x"5A",x"15",x"00",x"00",
																x"00",x"00",x"80",x"90",x"B8",x"58",x"8D",x"22",x"00",x"00",x"80",x"90",x"B8",x"58",x"8D",x"22",x"00",x"30",x"7B",x"6F",x"D5",x"AA",x"45",x"02",x"00",x"30",x"7B",x"6F",x"D5",x"AA",x"45",x"02",x"80",x"00",x"20",x"74",x"D0",x"A8",x"56",x"0A",x"80",x"00",x"20",x"74",x"D0",x"A8",x"56",x"0A",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"00",x"00",x"18",x"3C",x"3C",x"18",x"00",x"00",x"00",x"00",x"18",x"3C",x"3C",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"38",x"4C",x"C6",x"C6",x"C6",x"64",x"38",x"00",x"38",x"4C",x"C6",x"C6",x"C6",x"64",x"38",x"00",x"92",x"54",x"38",x"FF",x"38",x"54",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"C7",x"B3",x"39",x"39",x"39",x"9B",x"C7",x"FF",x"38",x"4C",x"C6",x"C6",x"C6",x"64",x"38",x"00",x"E7",x"C7",x"E7",x"E7",x"E7",x"E7",x"81",x"FF",x"18",x"38",x"18",x"18",x"18",x"18",x"7E",x"00",x"83",x"39",x"F1",x"C3",x"87",x"1F",x"01",x"FF",x"7C",x"C6",x"0E",x"3C",x"78",x"E0",x"FE",x"00",x"81",x"F3",x"E7",x"C3",x"F9",x"39",x"83",x"FF",x"7E",x"0C",x"18",x"3C",x"06",x"C6",x"7C",x"00",
																x"E3",x"C3",x"93",x"33",x"01",x"F3",x"F3",x"FF",x"1C",x"3C",x"6C",x"CC",x"FE",x"0C",x"0C",x"00",x"03",x"3F",x"03",x"F9",x"F9",x"39",x"83",x"FF",x"FC",x"C0",x"FC",x"06",x"06",x"C6",x"7C",x"00",x"C3",x"9F",x"3F",x"03",x"39",x"39",x"83",x"FF",x"3C",x"60",x"C0",x"FC",x"C6",x"C6",x"7C",x"00",x"01",x"39",x"F3",x"E7",x"CF",x"CF",x"CF",x"FF",x"FE",x"C6",x"0C",x"18",x"30",x"30",x"30",x"00",
																x"83",x"39",x"39",x"83",x"39",x"39",x"83",x"FF",x"7C",x"C6",x"C6",x"7C",x"C6",x"C6",x"7C",x"00",x"83",x"39",x"39",x"81",x"F9",x"F3",x"87",x"FF",x"7C",x"C6",x"C6",x"7E",x"06",x"0C",x"78",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"C6",x"C6",x"FC",x"C6",x"C6",x"FC",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3C",x"66",x"C0",x"C0",x"C0",x"66",x"3C",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"CC",x"C6",x"C6",x"C6",x"CC",x"F8",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"FE",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"C0",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3E",x"60",x"C0",x"CE",x"C6",x"66",x"3E",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1E",x"0C",x"0C",x"0C",x"0C",x"CC",x"78",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"CC",x"D8",x"F0",x"F8",x"DC",x"CE",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"C6",x"C6",x"C6",x"FC",x"C0",x"C0",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"38",x"6C",x"C6",x"C6",x"DE",x"6C",x"3A",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"C6",x"C6",x"FC",x"D8",x"CC",x"C6",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7C",x"C6",x"C0",x"7C",x"06",x"C6",x"7C",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"C6",x"6C",x"6C",x"38",x"38",x"10",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"C6",x"D6",x"FE",x"FE",x"EE",x"C6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"C6",x"6C",x"38",x"6C",x"C6",x"C6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"0E",x"1C",x"38",x"70",x"E0",x"FE",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7C",x"82",x"9A",x"A2",x"9A",x"82",x"7C",x"00",x"FF",x"BB",x"D7",x"EF",x"D7",x"BB",x"FF",x"FF",x"00",x"44",x"28",x"10",x"28",x"44",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7C",x"7C",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"E7",x"E7",x"FF",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",
																x"FF",x"FF",x"FF",x"03",x"03",x"FF",x"FF",x"FF",x"00",x"00",x"03",x"FF",x"FF",x"03",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"CD",x"CD",x"CD",x"CD",x"CD",x"F7",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"22",x"A2",x"AA",x"BE",x"BE",x"B6",x"22",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																x"FB",x"F3",x"F3",x"F3",x"F3",x"F3",x"FB",x"FF",x"04",x"0C",x"0C",x"0C",x"0C",x"0C",x"04",x"00",x"07",x"8B",x"F3",x"F3",x"F3",x"F3",x"CB",x"87",x"F8",x"74",x"0C",x"0C",x"0C",x"0C",x"34",x"78",x"7F",x"3F",x"3F",x"3F",x"3F",x"47",x"83",x"FF",x"80",x"C0",x"C0",x"C0",x"C0",x"B8",x"7C",x"00",x"FB",x"F3",x"F3",x"F3",x"F3",x"8B",x"07",x"FF",x"04",x"0C",x"0C",x"0C",x"0C",x"74",x"F8",x"00",
																x"7B",x"33",x"33",x"33",x"33",x"33",x"4B",x"87",x"84",x"CC",x"CC",x"CC",x"CC",x"CC",x"B4",x"78",x"83",x"47",x"3F",x"3F",x"3F",x"3F",x"4F",x"87",x"7C",x"B8",x"C0",x"C0",x"C0",x"C0",x"B0",x"78",x"7B",x"33",x"33",x"33",x"33",x"4B",x"87",x"FF",x"84",x"CC",x"CC",x"CC",x"CC",x"B4",x"78",x"00",x"07",x"8B",x"F3",x"F3",x"F3",x"F3",x"FB",x"FF",x"F8",x"74",x"0C",x"0C",x"0C",x"0C",x"04",x"00",
																x"87",x"4B",x"33",x"33",x"33",x"33",x"4B",x"87",x"78",x"B4",x"CC",x"CC",x"CC",x"CC",x"B4",x"78",x"87",x"4B",x"33",x"33",x"33",x"33",x"7B",x"FF",x"78",x"B4",x"CC",x"CC",x"CC",x"CC",x"84",x"00",x"FB",x"F3",x"F3",x"F3",x"F3",x"F3",x"FB",x"FF",x"04",x"0C",x"0C",x"0C",x"0C",x"0C",x"04",x"00",x"39",x"19",x"09",x"01",x"21",x"31",x"39",x"FF",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"00",
																x"FF",x"FF",x"C3",x"99",x"99",x"99",x"C3",x"FF",x"00",x"00",x"3C",x"66",x"66",x"66",x"3C",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"C0",x"D0",x"D0",x"E6",x"F7",x"D5",x"D5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"C2",x"C4",x"48",x"50",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"01",x"02",x"04",x"08",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"20",x"58",x"98",x"1E",x"1A",x"1A",x"1A",x"00",x"FF",x"FD",x"F9",x"F1",x"F1",x"D1",x"91",x"13",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"17",x"1F",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FD",x"F9",x"F1",x"F1",x"F1",x"F1",x"F3",x"00",x"00",x"00",x"00",x"00",x"20",x"60",x"E0",
																x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"02",x"06",x"0E",x"0E",x"2E",x"6E",x"EC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E8",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"11",x"11",x"11",x"11",x"11",x"11",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"F1",x"F1",x"F1",x"F1",x"F1",x"F1",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EE",x"EE",x"EE",x"EE",x"EE",x"EE",x"00",x"00",x"11",x"11",x"11",x"11",x"11",x"11",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"11",x"11",x"11",x"11",x"11",x"11",x"FF",x"FF",x"EE",x"EE",x"EE",x"EE",x"EE",x"EE",x"00",x"00",
																x"FF",x"80",x"C0",x"E0",x"F0",x"FF",x"FF",x"FF",x"00",x"7F",x"3F",x"1F",x"0F",x"00",x"00",x"00",x"FF",x"03",x"07",x"0F",x"1F",x"FF",x"FF",x"FF",x"00",x"FC",x"F8",x"F0",x"E0",x"00",x"00",x"00",x"FF",x"FF",x"F0",x"E0",x"C0",x"80",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"1F",x"0F",x"07",x"03",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"FF",x"80",x"C0",x"E0",x"F0",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"03",x"07",x"0F",x"1F",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F0",x"E0",x"C0",x"80",x"FF",x"FF",x"00",x"00",x"0F",x"1F",x"3F",x"7F",x"00",x"00",x"FF",x"FF",x"1F",x"0F",x"07",x"03",x"FF",x"FF",x"00",x"00",x"E0",x"F0",x"F8",x"FC",x"00",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"C0",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																x"3E",x"60",x"C0",x"CE",x"C6",x"66",x"3E",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E2",x"C0",x"80",x"E0",x"F2",x"FC",x"FF",x"00",x"1D",x"3F",x"7F",x"1F",x"0D",x"03",x"00",x"8F",x"17",x"0B",x"27",x"9F",x"2B",x"DF",x"FF",x"70",x"E8",x"F4",x"D8",x"60",x"D4",x"20",x"00",
																x"FF",x"FF",x"FC",x"E0",x"C0",x"F8",x"FE",x"FF",x"00",x"00",x"03",x"1F",x"3F",x"07",x"01",x"00",x"FF",x"F1",x"40",x"00",x"00",x"22",x"19",x"FC",x"00",x"0E",x"BF",x"FF",x"FF",x"DD",x"E6",x"03",x"88",x"00",x"05",x"02",x"94",x"4B",x"07",x"7F",x"77",x"FF",x"FA",x"FD",x"6B",x"B4",x"F8",x"80",x"FF",x"3F",x"47",x"0F",x"FF",x"7D",x"CF",x"E7",x"00",x"C0",x"B8",x"F0",x"00",x"82",x"30",x"18",
																x"00",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"00",x"08",x"08",x"00",x"08",x"08",x"00",x"00",x"08",x"08",x"08",x"00",x"08",x"08",x"00",x"00",x"08",x"08",
																x"08",x"00",x"08",x"08",x"08",x"00",x"00",x"08",x"08",x"00",x"08",x"08",x"08",x"00",x"00",x"08",x"08",x"08",x"00",x"08",x"08",x"08",x"00",x"00",x"08",x"08",x"00",x"08",x"08",x"08",x"00",x"00",x"00",x"08",x"08",x"00",x"08",x"08",x"08",x"00",x"00",x"08",x"08",x"00",x"08",x"08",x"08",x"00",x"00",x"08",x"08",x"00",x"00",x"08",x"08",x"08",x"00",x"08",x"08",x"00",x"00",x"08",x"08",x"08",
																x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",
																x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",
																x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"00",
																x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",
																x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",
																x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",
																x"1C",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",
																x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"1C",x"1C",x"1C",x"1C",x"1C",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",
																x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",
																x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",
																x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",
																x"FF",x"80",x"2F",x"40",x"00",x"00",x"80",x"FF",x"00",x"00",x"2F",x"40",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"01",x"F0",x"00",x"00",x"00",x"01",x"FF",x"00",x"00",x"F0",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",
																x"00",x"FD",x"FA",x"F4",x"E8",x"D0",x"90",x"20",x"00",x"03",x"06",x"0C",x"18",x"30",x"70",x"E0",x"FE",x"FC",x"F9",x"F2",x"E2",x"C4",x"88",x"10",x"01",x"03",x"07",x"0E",x"1E",x"3C",x"78",x"F0",x"40",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FC",x"F8",x"F0",x"E1",x"C2",x"84",x"08",x"01",x"03",x"07",x"0F",x"1F",x"3E",x"7C",x"F8",
																x"20",x"40",x"40",x"80",x"00",x"00",x"00",x"00",x"E0",x"C0",x"C0",x"80",x"00",x"00",x"00",x"00",x"FE",x"FC",x"F8",x"F0",x"E0",x"C1",x"81",x"02",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FE",x"08",x"10",x"20",x"40",x"80",x"00",x"00",x"00",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"01",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",
																x"04",x"08",x"10",x"20",x"20",x"40",x"80",x"00",x"FC",x"F8",x"F0",x"E0",x"E0",x"C0",x"80",x"00",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"02",x"04",x"04",x"08",x"10",x"20",x"40",x"80",x"FE",x"FC",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"01",x"02",x"04",x"08",x"10",x"10",x"20",x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"F0",x"E0",
																x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"04",x"08",x"10",x"FF",x"FF",x"FF",x"FE",x"FE",x"FC",x"F8",x"F0",x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"08",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"02",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",
																x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"BF",x"5F",x"2F",x"17",x"0B",x"09",x"04",x"00",x"C0",x"60",x"30",x"18",x"0C",x"0E",x"07",x"7F",x"3F",x"9F",x"4F",x"47",x"23",x"11",x"08",x"80",x"C0",x"E0",x"70",x"78",x"3C",x"1E",x"0F",x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",
																x"7F",x"3F",x"1F",x"0F",x"87",x"43",x"21",x"10",x"80",x"C0",x"E0",x"F0",x"F8",x"7C",x"3E",x"1F",x"04",x"02",x"02",x"01",x"00",x"00",x"00",x"00",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"7F",x"3F",x"1F",x"0F",x"07",x"83",x"81",x"40",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"7F",x"10",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"1F",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",
																x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"80",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"20",x"10",x"08",x"04",x"04",x"02",x"01",x"00",x"3F",x"1F",x"0F",x"07",x"07",x"03",x"01",x"00",x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"40",x"20",x"20",x"10",x"08",x"04",x"02",x"01",x"7F",x"3F",x"3F",x"1F",x"0F",x"07",x"03",x"01",
																x"00",x"80",x"40",x"20",x"10",x"08",x"08",x"04",x"FF",x"FF",x"7F",x"3F",x"1F",x"0F",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"40",x"20",x"10",x"08",x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"1F",x"0F",x"00",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",
																x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"40",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"18",x"18",x"FF",x"FF",x"FF",x"00",x"00",x"18",x"FF",x"FF",x"18",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",
																x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"CF",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"03",x"01",x"00",x"00",x"00",x"00",x"01",x"03",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"01",x"87",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"FE",x"78",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"83",x"01",x"38",x"00",x"00",x"00",x"00",x"00",x"7C",x"FE",x"C7",
																x"FF",x"FF",x"FF",x"FC",x"F0",x"E1",x"C7",x"CF",x"00",x"00",x"00",x"03",x"0F",x"1E",x"38",x"30",x"FF",x"FF",x"FF",x"3F",x"1F",x"8F",x"CF",x"CF",x"00",x"00",x"00",x"C0",x"E0",x"70",x"30",x"30",x"FF",x"C7",x"E1",x"F0",x"FC",x"FF",x"FF",x"FF",x"30",x"38",x"1E",x"0F",x"03",x"00",x"00",x"00",x"FF",x"CF",x"8F",x"1F",x"3F",x"FF",x"FF",x"FF",x"30",x"30",x"70",x"E0",x"C0",x"00",x"00",x"00",
																x"7F",x"3F",x"1F",x"8F",x"C7",x"E3",x"F1",x"F8",x"80",x"C0",x"E0",x"70",x"38",x"1C",x"0E",x"07",x"F8",x"F1",x"E3",x"C7",x"8F",x"1F",x"3F",x"7F",x"07",x"0E",x"1C",x"38",x"70",x"E0",x"C0",x"80",x"78",x"31",x"63",x"C7",x"8F",x"1B",x"31",x"78",x"87",x"CE",x"9C",x"38",x"70",x"E4",x"CE",x"87",x"CF",x"CF",x"FF",x"00",x"00",x"FF",x"CF",x"CF",x"30",x"30",x"00",x"FF",x"FF",x"00",x"30",x"30",
																x"F0",x"C0",x"87",x"1F",x"3F",x"3F",x"7F",x"7F",x"0F",x"3F",x"78",x"E0",x"C0",x"C0",x"80",x"80",x"1F",x"07",x"C3",x"F1",x"F9",x"F8",x"FC",x"FC",x"E0",x"F8",x"3C",x"0E",x"06",x"07",x"03",x"03",x"F8",x"F9",x"F1",x"F3",x"E3",x"87",x"0F",x"3F",x"07",x"06",x"0E",x"0C",x"1C",x"78",x"F0",x"C0",x"7F",x"1F",x"07",x"C0",x"F0",x"FF",x"FF",x"FF",x"80",x"E0",x"F8",x"3F",x"0F",x"00",x"00",x"00",
																x"F8",x"E1",x"83",x"0F",x"3F",x"FF",x"FF",x"FF",x"07",x"1E",x"7C",x"F0",x"C0",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"F8",x"E0",x"83",x"0F",x"3F",x"00",x"00",x"00",x"07",x"1F",x"7C",x"F0",x"C0",x"FF",x"FF",x"FF",x"3F",x"0F",x"83",x"E1",x"F8",x"00",x"00",x"00",x"C0",x"F0",x"7C",x"1E",x"07",x"F8",x"F0",x"E3",x"E7",x"C7",x"CF",x"CF",x"CF",x"07",x"0F",x"1C",x"18",x"38",x"30",x"30",x"30",
																x"F8",x"F1",x"E3",x"E7",x"C7",x"CF",x"CF",x"CF",x"07",x"0E",x"1C",x"18",x"38",x"30",x"30",x"30",x"7F",x"3F",x"3F",x"1F",x"9F",x"8F",x"CF",x"CF",x"80",x"C0",x"C0",x"E0",x"60",x"70",x"30",x"30",x"FF",x"CF",x"C7",x"E3",x"E3",x"F1",x"F8",x"FC",x"30",x"30",x"38",x"1C",x"1C",x"0E",x"07",x"03",x"FF",x"CF",x"8F",x"9F",x"9F",x"1F",x"3F",x"7F",x"30",x"30",x"70",x"60",x"60",x"E0",x"C0",x"80",
																x"CF",x"CF",x"8F",x"1F",x"3F",x"FE",x"FE",x"FC",x"30",x"30",x"70",x"E0",x"C0",x"01",x"01",x"03",x"7E",x"3E",x"3F",x"1F",x"9F",x"8F",x"CF",x"CF",x"81",x"C1",x"C0",x"E0",x"60",x"70",x"30",x"30",x"7C",x"3E",x"3F",x"1F",x"9F",x"8F",x"CF",x"CF",x"83",x"C1",x"C0",x"E0",x"60",x"70",x"30",x"30",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"03",x"0F",x"3F",x"7F",x"FF",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"07",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"03",x"03",x"37",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F9",x"FF",x"00",x"00",x"C0",x"F0",x"FC",x"F7",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"EF",x"00",x"00",x"00",x"00",x"C0",x"F0",x"DC",x"EE",
																x"FF",x"FF",x"FF",x"DF",x"FB",x"FD",x"FF",x"FF",x"C0",x"F8",x"FE",x"DF",x"FB",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"FF",x"00",x"00",x"F0",x"FC",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"E0",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"01",x"03",x"0F",x"1F",x"7F",x"FF",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"03",x"07",x"0F",x"1F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"03",x"07",x"07",x"0F",x"1F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"DF",x"EF",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F3",x"FF",x"FF",x"C0",x"E0",x"F8",x"EF",x"F7",x"F3",x"FF",x"FF",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"FC",
																x"FF",x"FF",x"FF",x"BF",x"DF",x"F7",x"FF",x"FF",x"00",x"80",x"C0",x"A0",x"D8",x"F4",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"66",x"66",x"67",x"66",x"66",x"F6",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E1",x"33",x"36",x"E6",x"C6",x"63",x"31",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E6",x"36",x"06",x"06",x"06",x"36",x"E3",x"00",
																x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"37",x"33",x"33",x"33",x"33",x"33",x"E7",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"0C",x"0C",x"0C",x"0C",x"0C",x"8C",x"00",x"FF",x"FC",x"F0",x"E0",x"C0",x"C0",x"80",x"80",x"00",x"03",x"0F",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF",x"3F",x"0F",x"07",x"03",x"03",x"01",x"01",x"00",x"C0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",
																x"80",x"80",x"C0",x"C0",x"E0",x"F0",x"FC",x"FF",x"7F",x"7F",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"01",x"01",x"03",x"03",x"07",x"0F",x"3F",x"FF",x"FE",x"FE",x"FC",x"FC",x"F8",x"F0",x"C0",x"00",x"00",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01");
	
	constant KUNG_FU_CHR_ROM : CHR_ROM_ARRAY := (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"A0",x"A0",x"A0",x"A0",x"A0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4E",x"CA",x"4A",x"4A",x"4A",x"4A",x"4E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EE",x"2A",x"2A",x"4A",x"8A",x"8A",x"EE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EE",x"AA",x"2A",x"6A",x"2A",x"AA",x"EE",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2E",x"6A",x"AA",x"AA",x"AA",x"FA",x"2E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EE",x"8A",x"8A",x"EA",x"2A",x"AA",x"EE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EE",x"AA",x"8A",x"EA",x"AA",x"AA",x"EE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EE",x"AA",x"AA",x"EA",x"AA",x"AA",x"EE",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EE",x"AA",x"AA",x"AA",x"AA",x"AA",x"EE",x"00",x"00",x"20",x"40",x"40",x"20",x"00",x"00",x"00",x"66",x"DF",x"BF",x"BF",x"DF",x"7E",x"3C",x"18",x"00",x"00",x"04",x"07",x"07",x"04",x"00",x"00",x"00",x"00",x"04",x"FC",x"7C",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"4A",x"2C",x"3E",x"78",x"3C",x"56",x"81",
																	x"3E",x"7F",x"77",x"C3",x"81",x"00",x"00",x"00",x"3C",x"7E",x"66",x"C3",x"81",x"00",x"00",x"00",x"38",x"70",x"F0",x"E0",x"E0",x"E0",x"60",x"30",x"30",x"60",x"E0",x"C0",x"C0",x"E0",x"60",x"30",x"39",x"7C",x"CE",x"87",x"84",x"CF",x"7C",x"3A",x"00",x"00",x"30",x"78",x"78",x"30",x"00",x"00",x"3E",x"78",x"FF",x"CE",x"CF",x"FE",x"7C",x"3D",x"00",x"00",x"00",x"30",x"30",x"00",x"00",x"00",
																	x"00",x"0B",x"1F",x"1F",x"1F",x"1F",x"0F",x"1F",x"00",x"0B",x"1F",x"1F",x"17",x"02",x"0A",x"00",x"0F",x"0F",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"03",x"0F",x"0F",x"0F",x"0F",x"0F",x"2F",x"AF",x"E7",x"E7",x"67",x"03",x"03",x"0F",x"0F",x"0F",x"1C",x"1E",x"18",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"1F",x"1F",x"3F",x"3F",
																	x"00",x"00",x"08",x"1C",x"FC",x"7C",x"3C",x"08",x"3F",x"1E",x"06",x"00",x"E0",x"7C",x"3C",x"08",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"40",x"40",x"80",x"80",x"00",x"C0",x"80",x"80",x"00",x"00",x"80",x"80",x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"80",x"80",x"C0",x"C0",x"80",x"80",x"80",x"90",x"FC",x"FC",x"FC",x"FC",x"FC",x"78",x"78",x"70",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F8",x"F0",x"F8",x"F8",x"D8",x"BC",x"7C",x"00",x"00",x"00",x"0E",x"0F",x"07",x"0E",x"3C",x"7E",x"3E",x"3E",x"30",x"11",x"03",x"0E",x"3C",x"00",x"02",x"07",x"07",x"07",x"07",x"03",x"07",x"00",x"02",x"07",x"07",x"05",x"00",x"02",x"00",x"00",x"03",x"01",x"01",x"03",x"03",x"07",x"07",x"00",x"00",x"00",x"00",x"03",x"03",x"07",x"07",
																	x"07",x"07",x"07",x"07",x"03",x"03",x"03",x"03",x"07",x"07",x"07",x"07",x"03",x"03",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0F",x"07",x"07",x"03",x"03",x"00",x"03",x"07",x"30",x"F8",x"F8",x"F0",x"C0",x"E0",x"E0",x"E0",x"00",x"80",x"80",x"CC",x"FC",x"BC",x"9C",x"1E",
																	x"E0",x"E0",x"C0",x"C0",x"00",x"04",x"04",x"0C",x"3E",x"3E",x"3E",x"FC",x"FC",x"FC",x"FC",x"FC",x"9C",x"FC",x"FC",x"F8",x"F8",x"F8",x"F8",x"FC",x"FC",x"FC",x"FC",x"F8",x"F8",x"F8",x"F8",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F0",x"E0",x"C0",x"80",x"C0",x"00",x"10",x"10",x"30",x"F0",x"E0",x"E0",x"C0",x"E0",x"F0",x"F0",x"D0",x"30",x"20",x"E0",x"C0",
																	x"3F",x"9B",x"F8",x"30",x"F0",x"20",x"60",x"07",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"C0",x"E0",x"E0",x"E0",x"C0",x"40",x"00",x"E0",x"00",x"00",x"00",x"38",x"2A",x"7E",x"3C",x"0C",x"18",x"3E",x"7C",x"07",x"14",x"01",x"02",x"00",x"06",x"0F",x"0F",x"07",x"C1",x"E0",x"E1",x"07",x"1E",x"3F",x"3F",x"3F",x"7F",x"3F",x"3E",x"1E",
																	x"1E",x"3D",x"7B",x"77",x"73",x"71",x"30",x"00",x"1E",x"3F",x"7F",x"77",x"73",x"71",x"00",x"F1",x"00",x"00",x"80",x"80",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"80",x"80",x"C0",x"C0",x"00",x"00",x"C0",x"00",x"00",x"80",x"C0",x"C0",x"80",x"00",x"00",x"00",x"00",x"80",x"C0",x"A0",x"40",x"80",x"06",x"0E",x"0E",x"0E",x"1C",x"3C",x"78",x"66",x"1E",x"3E",x"3E",x"3E",x"3E",x"1E",x"1E",x"1E",
																	x"3E",x"3C",x"38",x"3C",x"1C",x"1C",x"0C",x"00",x"3E",x"3C",x"38",x"3C",x"1C",x"08",x"32",x"1C",x"00",x"02",x"0F",x"0F",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"18",x"3C",x"FC",x"F8",x"E0",x"00",x"00",x"06",x"1E",x"3F",x"FF",x"FF",x"FF",x"1F",x"1F",x"1E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"0F",x"1F",x"1F",x"3F",
																	x"07",x"03",x"1B",x"0D",x"3D",x"2D",x"08",x"00",x"3F",x"7F",x"E7",x"F3",x"C3",x"D1",x"40",x"00",x"00",x"00",x"00",x"00",x"20",x"70",x"70",x"70",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",x"F0",x"6C",x"5C",x"FC",x"F8",x"F0",x"E0",x"C0",x"00",x"EA",x"DA",x"FA",x"FE",x"F2",x"E0",x"C0",x"00",x"00",x"00",x"00",x"1E",x"3E",x"3E",x"3D",x"3B",x"00",x"00",x"18",x"2E",x"5E",x"5E",x"3D",x"3F",
																	x"7B",x"47",x"0F",x"07",x"03",x"00",x"00",x"00",x"7F",x"7F",x"7F",x"7F",x"7F",x"3F",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"E0",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"B8",x"70",x"78",x"D8",x"10",x"00",x"00",x"00",x"80",x"88",x"84",x"A4",x"EC",x"FC",x"38",x"00",x"00",x"00",x"00",x"03",x"01",x"07",x"03",x"0F",x"00",x"03",x"07",x"00",x"02",x"00",x"01",x"0F",
																	x"1F",x"0C",x"03",x"0F",x"1F",x"1F",x"0E",x"00",x"1F",x"0F",x"03",x"0F",x"1F",x"1F",x"10",x"3C",x"00",x"00",x"00",x"00",x"40",x"80",x"C0",x"E0",x"00",x"C0",x"E0",x"E0",x"B0",x"70",x"F8",x"FC",x"C0",x"00",x"E0",x"F0",x"F8",x"F8",x"F0",x"E0",x"FE",x"FE",x"FE",x"FE",x"FC",x"F8",x"F0",x"E0",x"00",x"0F",x"1F",x"00",x"03",x"0F",x"0F",x"1F",x"00",x"0F",x"1F",x"1F",x"1F",x"02",x"08",x"00",
																	x"00",x"00",x"80",x"00",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"50",x"40",x"00",x"07",x"0F",x"00",x"01",x"07",x"07",x"0F",x"00",x"07",x"0F",x"0F",x"0F",x"01",x"04",x"00",x"07",x"07",x"03",x"03",x"07",x"07",x"0F",x"0F",x"00",x"00",x"00",x"01",x"07",x"07",x"0F",x"0F",x"2F",x"EF",x"60",x"60",x"60",x"00",x"00",x"03",x"0F",x"0F",x"1F",x"1F",x"1F",x"0F",x"03",x"03",
																	x"00",x"00",x"00",x"20",x"30",x"38",x"7C",x"78",x"00",x"03",x"07",x"2E",x"1C",x"08",x"04",x"00",x"30",x"80",x"E0",x"00",x"E0",x"E0",x"E0",x"E0",x"40",x"F0",x"F0",x"F0",x"F0",x"70",x"28",x"20",x"C0",x"C0",x"80",x"E0",x"80",x"80",x"00",x"00",x"60",x"70",x"70",x"F0",x"E0",x"F0",x"F0",x"F8",x"00",x"00",x"00",x"08",x"08",x"18",x"38",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",
																	x"00",x"00",x"20",x"E0",x"60",x"60",x"20",x"00",x"00",x"00",x"00",x"1E",x"1F",x"1F",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"3C",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"7E",x"7F",x"0F",x"3F",x"3F",x"7F",x"3F",x"3E",x"0E",x"0E",x"7F",x"0B",x"21",x"03",x"C3",x"C1",x"F3",x"F7",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"FF",x"7F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"1F",x"3F",x"7F",x"FF",x"FE",x"FE",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"40",x"00",x"E0",x"F0",x"F8",x"F8",x"00",x"80",x"C0",x"E0",x"C0",x"C0",x"80",x"E0",x"FC",x"FC",x"FE",x"FE",x"FE",x"FC",x"FC",x"98",x"F0",x"70",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"88",x"98",x"F0",x"F0",x"F8",x"FC",x"FE",
																	x"00",x"00",x"02",x"07",x"0F",x"07",x"0E",x"1C",x"FE",x"FE",x"7C",x"39",x"11",x"03",x"0E",x"1C",x"00",x"80",x"C0",x"00",x"E0",x"E0",x"E0",x"E0",x"00",x"80",x"C0",x"E0",x"F0",x"70",x"28",x"20",x"C0",x"C0",x"80",x"C0",x"90",x"80",x"00",x"00",x"40",x"40",x"00",x"C0",x"F0",x"F0",x"F8",x"F8",x"00",x"08",x"08",x"08",x"08",x"19",x"38",x"F8",x"F8",x"FC",x"FF",x"FF",x"FF",x"FE",x"F8",x"F8",
																	x"00",x"00",x"00",x"50",x"F0",x"F0",x"70",x"00",x"00",x"00",x"00",x"90",x"3E",x"1F",x"10",x"00",x"0F",x"3F",x"3F",x"7F",x"3F",x"3E",x"0F",x"0F",x"7F",x"0B",x"21",x"03",x"03",x"01",x"03",x"07",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"3F",x"7F",x"FF",x"FF",x"00",x"00",x"08",x"1C",x"3C",x"1C",x"08",x"00",x"01",x"03",x"07",x"03",x"03",x"03",x"02",x"00",
																	x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"EF",x"DF",x"BF",x"7F",x"FF",x"FE",x"FC",x"0C",x"06",x"03",x"03",x"37",x"3F",x"7E",x"78",x"0C",x"06",x"03",x"03",x"17",x"0E",x"04",x"00",x"0C",x"1E",x"FF",x"F7",x"E3",x"C3",x"06",x"0C",x"0C",x"1E",x"33",x"11",x"01",x"03",x"06",x"0C",x"00",x"00",x"F8",x"6C",x"3C",x"0E",x"1E",x"7E",x"00",x"00",x"E0",x"74",x"BC",x"7E",x"1E",x"7E",
																	x"0E",x"1C",x"38",x"70",x"79",x"79",x"3F",x"1F",x"06",x"04",x"08",x"10",x"19",x"0F",x"07",x"01",x"00",x"00",x"00",x"00",x"C0",x"C0",x"E8",x"3D",x"00",x"00",x"00",x"00",x"E0",x"F0",x"F8",x"3F",x"00",x"00",x"40",x"80",x"C8",x"F8",x"98",x"0E",x"00",x"00",x"60",x"F0",x"F8",x"F8",x"9C",x"0E",x"01",x"01",x"07",x"05",x"01",x"00",x"01",x"03",x"01",x"03",x"07",x"01",x"00",x"00",x"02",x"03",
																	x"0E",x"9E",x"7C",x"78",x"F8",x"78",x"F0",x"70",x"02",x"87",x"4F",x"58",x"DC",x"7E",x"D8",x"1C",x"78",x"F8",x"FC",x"7C",x"3C",x"BC",x"7C",x"FC",x"18",x"9E",x"8C",x"4F",x"0E",x"8C",x"4F",x"DE",x"78",x"F0",x"F0",x"70",x"78",x"3C",x"1F",x"0F",x"78",x"9C",x"B8",x"30",x"1C",x"0E",x"07",x"01",x"00",x"14",x"18",x"24",x"70",x"C0",x"C0",x"80",x"15",x"2A",x"3F",x"7A",x"6C",x"F0",x"C0",x"80",
																	x"0F",x"1F",x"3F",x"3F",x"5F",x"CB",x"DF",x"DF",x"0F",x"1F",x"3F",x"31",x"44",x"CD",x"C1",x"C0",x"CF",x"CF",x"C7",x"C7",x"CF",x"CF",x"CF",x"CF",x"C0",x"C0",x"C0",x"C3",x"CF",x"CF",x"CF",x"CF",x"80",x"00",x"E0",x"C0",x"80",x"00",x"00",x"00",x"80",x"00",x"E0",x"F0",x"F8",x"F8",x"FC",x"FC",x"0F",x"1F",x"3F",x"3F",x"1F",x"0B",x"1F",x"1F",x"0F",x"1F",x"3F",x"31",x"04",x"0D",x"01",x"00",
																	x"06",x"0E",x"8C",x"DC",x"F8",x"F8",x"F8",x"F8",x"06",x"0E",x"8C",x"DC",x"D8",x"C8",x"40",x"40",x"80",x"40",x"E0",x"F0",x"80",x"00",x"00",x"00",x"F8",x"F8",x"F0",x"F0",x"F0",x"F8",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"30",x"70",x"60",x"C0",x"C0",x"80",x"80",x"00",x"30",x"70",x"60",x"C0",x"C0",x"80",x"80",x"00",
																	x"80",x"F0",x"F0",x"78",x"70",x"30",x"00",x"00",x"80",x"C0",x"E0",x"26",x"0F",x"0F",x"1F",x"07",x"00",x"00",x"00",x"00",x"3C",x"7C",x"FE",x"FF",x"00",x"00",x"00",x"00",x"3C",x"7C",x"FE",x"C7",x"7F",x"2F",x"7F",x"7F",x"0E",x"3F",x"2F",x"0F",x"13",x"37",x"05",x"01",x"B2",x"C3",x"DF",x"FF",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"F0",x"F8",x"F8",
																	x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"70",x"38",x"1C",x"0E",x"07",x"80",x"C0",x"E0",x"70",x"38",x"1C",x"0E",x"07",x"00",x"00",x"00",x"07",x"0F",x"1F",x"1F",x"0F",x"00",x"00",x"00",x"07",x"0F",x"1F",x"18",x"02",x"05",x"0F",x"0F",x"07",x"07",x"03",x"03",x"07",x"1E",x"30",x"30",x"38",x"38",x"1D",x"0F",x"00",
																	x"07",x"07",x"03",x"01",x"01",x"01",x"00",x"00",x"08",x"38",x"7C",x"7E",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"10",x"3C",x"3C",x"78",x"F0",x"FC",x"7C",x"78",x"28",x"04",x"0C",x"78",x"F0",x"06",x"0E",x"0C",x"9C",x"F8",x"F8",x"F8",x"F8",x"06",x"0E",x"0C",x"9C",x"98",x"C8",x"E0",x"60",x"E0",x"E0",x"E0",x"DC",x"E6",x"C3",x"81",x"81",x"E0",x"A0",x"20",x"5C",x"7E",x"FF",x"FF",x"FF",
																	x"81",x"81",x"01",x"01",x"03",x"C6",x"FC",x"00",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"3F",x"3F",x"1F",x"1F",x"0F",x"0F",x"06",x"20",x"30",x"70",x"78",x"38",x"38",x"18",x"38",x"20",x"30",x"90",x"98",x"C8",x"88",x"08",x"38",x"00",x"00",x"00",x"00",x"3C",x"FC",x"FC",x"18",x"00",x"00",x"00",x"01",x"03",x"F3",x"E3",x"03",
																	x"00",x"00",x"00",x"0F",x"1F",x"3F",x"3F",x"1F",x"00",x"00",x"00",x"0F",x"1F",x"3F",x"31",x"04",x"0B",x"1F",x"1F",x"03",x"0F",x"0F",x"07",x"07",x"0D",x"01",x"00",x"EC",x"F0",x"F5",x"FF",x"F8",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"B0",x"FC",x"E6",x"C2",x"82",x"C0",x"40",x"40",x"30",x"FC",x"FE",x"FE",x"FE",
																	x"00",x"00",x"00",x"00",x"00",x"FF",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"7F",x"00",x"00",x"3C",x"7A",x"FD",x"FD",x"5F",x"FF",x"BF",x"00",x"00",x"04",x"02",x"02",x"10",x"00",x"00",x"7F",x"7F",x"7F",x"1F",x"1F",x"1F",x"1F",x"1F",x"01",x"03",x"06",x"04",x"0C",x"1C",x"1C",x"1E",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"7F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"1F",
																	x"FF",x"DF",x"EE",x"E0",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"1F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"00",x"E0",x"F0",x"D8",x"EC",x"F4",x"F6",x"FE",x"80",x"00",x"00",x"20",x"10",x"08",x"08",x"00",x"FF",x"EF",x"F7",x"F7",x"F7",x"FE",x"FE",x"FE",x"00",x"90",x"C8",x"E8",x"E8",x"E0",x"E0",x"E0",
																	x"FE",x"BC",x"3E",x"1E",x"0C",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"E0",x"F2",x"FC",x"FC",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"E8",x"D8",x"B8",x"7C",x"FC",x"7E",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"1F",x"3F",x"3F",x"3F",x"3F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F0",x"F0",x"E0",x"E0",x"E0",
																	x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"7F",x"3F",x"3F",x"33",x"21",x"20",x"20",x"30",x"1E",x"FF",x"FF",x"FF",x"FF",x"F7",x"8F",x"FF",x"FE",x"00",x"80",x"C0",x"E0",x"08",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"3C",x"7E",x"FE",x"3F",x"3F",x"3E",x"1E",x"04",x"00",x"42",x"FE",x"FE",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"F8",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F8",x"FC",x"FC",x"7E",x"7E",x"00",x"00",x"00",x"0C",x"0E",x"0F",x"3F",x"7F",x"7E",x"7F",x"3F",x"33",x"10",x"01",x"31",x"7F",x"00",x"38",x"4F",x"BF",x"FF",x"EF",x"70",x"00",x"00",x"00",x"30",x"40",x"00",x"00",x"00",x"00",x"00",x"1F",x"F1",x"DF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"0E",x"20",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"3C",x"7A",x"FD",x"FD",x"5F",x"FF",x"00",x"00",x"00",x"04",x"02",x"02",x"10",x"00",x"BF",x"FF",x"8F",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"F9",x"B2",x"E4",x"84",x"CC",x"FC",x"FE",x"7F",x"3F",x"3F",x"3F",x"3F",x"3F",x"1F",x"1F",x"7F",x"3F",x"3F",x"3F",x"3F",x"3F",x"1E",x"1E",x"0F",x"07",x"0F",x"0C",x"00",x"00",x"00",x"00",x"0C",x"04",x"0C",x"0F",x"0F",x"0F",x"0F",x"0F",
																	x"00",x"C0",x"E0",x"B8",x"CC",x"F6",x"FE",x"FF",x"00",x"00",x"00",x"40",x"30",x"08",x"00",x"00",x"FF",x"FF",x"FF",x"F7",x"F7",x"EE",x"FE",x"FC",x"C0",x"F0",x"F0",x"E8",x"E8",x"D0",x"40",x"00",x"FC",x"F8",x"E0",x"00",x"00",x"00",x"00",x"00",x"04",x"0E",x"1E",x"FE",x"FE",x"FC",x"FC",x"F8",x"FF",x"E3",x"C1",x"80",x"00",x"00",x"00",x"00",x"0F",x"1F",x"3F",x"7F",x"7F",x"7F",x"7F",x"7F",
																	x"00",x"00",x"98",x"FC",x"FC",x"7C",x"3C",x"18",x"7F",x"3F",x"86",x"C2",x"F0",x"7C",x"3C",x"18",x"40",x"60",x"70",x"78",x"7C",x"3C",x"3C",x"38",x"40",x"67",x"67",x"67",x"63",x"33",x"33",x"33",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"00",x"07",x"0F",x"1F",x"1F",x"0B",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",
																	x"17",x"0F",x"01",x"0F",x"EF",x"F7",x"D7",x"E7",x"00",x"0F",x"0E",x"0C",x"01",x"06",x"06",x"06",x"EF",x"FF",x"FF",x"7F",x"7F",x"3F",x"0F",x"0F",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"0F",x"7F",x"00",x"00",x"80",x"40",x"A0",x"A0",x"E0",x"E0",x"00",x"00",x"00",x"80",x"40",x"40",x"00",x"00",x"E0",x"E0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",x"00",x"20",x"40",x"80",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"01",x"00",x"01",x"03",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"E0",x"60",x"F0",x"FE",x"FF",x"00",x"F0",x"B8",x"18",x"98",x"0C",x"1E",x"3F",x"7F",x"C7",x"83",x"83",x"83",x"C1",x"C1",x"E0",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"E0",x"61",x"42",x"33",x"7B",x"FE",x"30",x"FF",x"FF",x"7F",x"7F",x"0F",x"47",x"D7",x"4F",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"1F",x"7F",x"7F",x"FE",x"FC",x"7E",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"F8",x"FF",x"FB",x"FB",x"79",x"7D",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"70",x"70",x"E0",x"C0",x"F0",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"02",x"06",x"0F",x"0E",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"05",x"0F",x"0F",x"07",
																	x"00",x"00",x"00",x"00",x"00",x"20",x"FE",x"3F",x"00",x"00",x"00",x"00",x"78",x"DC",x"1E",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"3F",x"C0",x"68",x"6C",x"FE",x"FC",x"78",x"28",x"00",x"0C",x"06",x"13",x"01",x"03",x"07",x"16",x"3C",x"00",x"00",x"00",x"00",x"03",x"00",x"03",x"07",x"00",x"00",x"01",x"03",x"00",x"01",x"00",x"00",
																	x"E0",x"60",x"60",x"41",x"01",x"01",x"01",x"00",x"10",x"19",x"1B",x"3F",x"3F",x"1F",x"0F",x"03",x"00",x"00",x"00",x"80",x"C0",x"C0",x"FC",x"FE",x"00",x"00",x"E0",x"70",x"30",x"30",x"1C",x"3E",x"FF",x"8F",x"87",x"07",x"03",x"01",x"81",x"E0",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
																	x"01",x"00",x"00",x"01",x"01",x"01",x"01",x"20",x"00",x"01",x"01",x"03",x"03",x"07",x"1F",x"1F",x"70",x"F0",x"30",x"10",x"00",x"00",x"00",x"00",x"0E",x"0C",x"08",x"00",x"00",x"00",x"00",x"00",x"30",x"D0",x"54",x"FC",x"F8",x"70",x"70",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"7E",x"7C",x"3C",x"18",x"20",x"10",x"0E",x"07",x"07",x"0F",x"0F",x"0F",x"27",x"17",x"0F",
																	x"03",x"01",x"03",x"03",x"0B",x"09",x"04",x"64",x"7F",x"FE",x"FC",x"FC",x"FC",x"FE",x"FF",x"1F",x"00",x"00",x"00",x"0C",x"1E",x"3E",x"7E",x"F0",x"01",x"03",x"07",x"03",x"01",x"02",x"7E",x"F0",x"70",x"78",x"78",x"70",x"60",x"E0",x"C0",x"00",x"88",x"88",x"98",x"B0",x"E0",x"E0",x"C0",x"00",x"04",x"2E",x"7F",x"3F",x"9F",x"DF",x"FF",x"3F",x"04",x"0E",x"03",x"0B",x"03",x"03",x"07",x"03",
																	x"7A",x"20",x"0E",x"1F",x"1F",x"1F",x"1F",x"1F",x"86",x"DE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FE",x"FE",x"FE",x"3C",x"80",x"00",x"00",x"F9",x"00",x"00",x"00",x"C0",x"60",x"C0",x"80",x"70",x"41",x"03",x"03",x"07",x"07",x"07",x"07",x"0F",x"3F",x"7F",x"3F",x"1F",x"07",x"07",x"07",x"FA",x"F8",x"F0",x"E0",x"E0",x"E0",x"E6",x"EE",x"82",x"DE",x"FE",x"FF",x"FF",x"FF",x"F9",x"F0",
																	x"0D",x"8F",x"79",x"EF",x"0F",x"DF",x"FE",x"8F",x"0E",x"9F",x"FF",x"FF",x"7F",x"BF",x"FB",x"83",x"60",x"80",x"C0",x"40",x"00",x"80",x"00",x"00",x"80",x"60",x"F0",x"C8",x"E0",x"90",x"C0",x"60",x"38",x"78",x"50",x"01",x"01",x"01",x"01",x"02",x"06",x"07",x"0F",x"0F",x"03",x"01",x"01",x"03",x"18",x"38",x"3C",x"3E",x"3F",x"1F",x"03",x"00",x"07",x"07",x"03",x"17",x"3F",x"3F",x"3F",x"7F",
																	x"3E",x"7F",x"9F",x"0F",x"0F",x"0F",x"0F",x"0F",x"3E",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1E",x"3E",x"7C",x"FC",x"38",x"C0",x"E0",x"F0",x"FE",x"FE",x"FC",x"FC",x"F8",x"E0",x"E0",x"F0",x"10",x"70",x"70",x"30",x"38",x"3C",x"1F",x"6C",x"00",x"00",x"00",x"20",x"38",x"3C",x"1F",x"6F",x"F0",x"FC",x"FC",x"FE",x"EF",x"6F",x"5F",x"1F",x"F3",x"FF",x"FF",x"FF",x"EF",x"0F",x"9F",x"DF",
																	x"3F",x"3C",x"38",x"38",x"18",x"08",x"00",x"00",x"BF",x"BC",x"38",x"34",x"14",x"04",x"04",x"04",x"00",x"18",x"2C",x"1A",x"0E",x"2C",x"3C",x"18",x"0C",x"06",x"13",x"05",x"01",x"03",x"C3",x"E6",x"00",x"18",x"3C",x"3A",x"72",x"BE",x"BE",x"BC",x"F8",x"F8",x"FC",x"F8",x"F0",x"F8",x"B8",x"BC",x"00",x"07",x"0F",x"3F",x"3B",x"3F",x"1F",x"0F",x"00",x"00",x"02",x"01",x"00",x"20",x"10",x"08",
																	x"80",x"C0",x"C0",x"E0",x"F0",x"F0",x"70",x"30",x"83",x"9F",x"BF",x"9F",x"CF",x"CF",x"6F",x"2F",x"0F",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"EF",x"5F",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"80",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F0",x"E0",x"C0",x"C0",x"80",x"80",x"00",
																	x"00",x"07",x"0F",x"1F",x"0F",x"07",x"17",x"3B",x"00",x"07",x"0F",x"1F",x"1E",x"1C",x"1C",x"38",x"79",x"70",x"7C",x"3E",x"DE",x"FC",x"FC",x"FF",x"7E",x"7F",x"73",x"21",x"C1",x"C3",x"FF",x"C7",x"F8",x"FE",x"C0",x"C0",x"80",x"87",x"C0",x"F0",x"F6",x"DE",x"FE",x"FF",x"FF",x"F8",x"FF",x"FF",x"FE",x"C0",x"C1",x"C3",x"43",x"C3",x"83",x"80",x"FF",x"C1",x"C0",x"C0",x"40",x"C0",x"80",x"87",
																	x"00",x"80",x"C0",x"E0",x"C0",x"C0",x"E0",x"C0",x"00",x"80",x"C0",x"60",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"9C",x"DC",x"7C",x"00",x"00",x"00",x"F8",x"FC",x"60",x"20",x"80",x"FC",x"DC",x"DC",x"DC",x"D6",x"D0",x"40",x"00",x"10",x"10",x"10",x"50",x"58",x"D7",x"C0",x"C0",
																	x"00",x"00",x"00",x"00",x"00",x"1C",x"3E",x"7F",x"00",x"00",x"00",x"00",x"00",x"1C",x"3E",x"7F",x"3F",x"3E",x"DE",x"FF",x"EE",x"F1",x"7B",x"7B",x"7B",x"F0",x"E4",x"E0",x"F0",x"E8",x"44",x"44",x"5E",x"5E",x"4C",x"00",x"00",x"00",x"00",x"00",x"21",x"21",x"32",x"3E",x"76",x"60",x"60",x"32",x"00",x"00",x"00",x"10",x"10",x"20",x"20",x"70",x"3C",x"1C",x"3C",x"28",x"68",x"10",x"10",x"00",
																	x"60",x"48",x"4C",x"1A",x"0B",x"0B",x"07",x"32",x"80",x"80",x"80",x"C0",x"B0",x"90",x"19",x"3E",x"00",x"00",x"03",x"07",x"0F",x"0F",x"1F",x"1E",x"00",x"00",x"00",x"00",x"0C",x"0E",x"07",x"03",x"1C",x"18",x"01",x"03",x"07",x"03",x"00",x"00",x"03",x"07",x"0E",x"0C",x"00",x"00",x"00",x"00",x"80",x"44",x"31",x"13",x"02",x"00",x"1A",x"30",x"07",x"0F",x"0F",x"0E",x"3D",x"7F",x"F5",x"EF",
																	x"00",x"00",x"10",x"00",x"00",x"00",x"02",x"00",x"02",x"10",x"28",x"10",x"06",x"8E",x"0C",x"01",x"00",x"00",x"0C",x"1F",x"3E",x"3C",x"00",x"00",x"60",x"10",x"00",x"09",x"19",x"01",x"02",x"0C",x"00",x"00",x"00",x"80",x"F0",x"BC",x"A7",x"68",x"00",x"00",x"00",x"80",x"F0",x"4C",x"5F",x"10",x"07",x"03",x"0D",x"1F",x"3E",x"3C",x"00",x"00",x"67",x"13",x"01",x"09",x"19",x"01",x"02",x"0C",
																	x"E0",x"6C",x"FE",x"BF",x"FF",x"B0",x"A0",x"68",x"E0",x"EC",x"F2",x"F3",x"FF",x"40",x"58",x"10",x"00",x"03",x"04",x"03",x"08",x"18",x"1C",x"0F",x"00",x"00",x"03",x"04",x"07",x"07",x"03",x"10",x"0F",x"0A",x"02",x"00",x"00",x"00",x"00",x"00",x"10",x"15",x"0D",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"1F",x"1F",x"00",x"00",x"02",x"01",x"06",x"09",x"09",x"16",
																	x"00",x"00",x"18",x"38",x"38",x"00",x"00",x"00",x"00",x"00",x"08",x"1C",x"34",x"18",x"00",x"00",x"00",x"12",x"0C",x"00",x"08",x"04",x"07",x"03",x"3F",x"3F",x"3F",x"1F",x"3F",x"7F",x"7F",x"3F",x"00",x"12",x"0C",x"00",x"00",x"02",x"01",x"00",x"1F",x"1F",x"0F",x"1F",x"1F",x"0F",x"07",x"01",x"00",x"00",x"40",x"20",x"08",x"46",x"23",x"42",x"04",x"00",x"42",x"28",x"1C",x"5E",x"2F",x"F3",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"09",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"04",x"03",x"0F",x"CF",x"EF",x"EF",x"E7",x"E7",x"67",x"03",x"03",x"CF",x"CF",x"4F",x"1C",x"1E",x"18",x"04",x"04",x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"03",x"03",x"01",x"01",x"00",x"00",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"00",x"C0",x"E0",x"80",x"00",x"00",x"C0",x"C0",x"80",x"C0",x"E0",x"80",x"00",x"00",x"00",x"00",x"00",x"3C",x"76",x"7F",x"3F",x"1F",x"00",x"00",x"00",x"30",x"7A",x"7F",x"27",x"17",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"30",x"02",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"D8",x"70",x"E0",x"20",x"80",x"00",x"00",x"00",x"70",x"A8",x"10",x"F0",x"60",x"C0",x"00",x"00",x"00",x"00",x"04",x"02",x"00",x"08",x"06",x"00",x"03",x"0F",x"1F",x"1F",x"0F",x"1F",x"3F",x"3F",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"BD",x"66",x"5E",x"5E",x"66",x"BD",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E7",x"C3",x"C3",x"E7",x"E7",x"FF",x"E7",x"FF",x"00",x"00",x"00",x"00",x"00",x"08",x"A4",x"FE",x"00",x"00",x"00",x"60",x"A8",x"F4",x"5A",x"01",x"00",x"00",x"00",x"00",x"34",x"1E",x"AD",x"FF",x"40",x"E2",x"34",x"FE",x"CB",x"E1",x"52",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"05",x"03",x"0F",x"00",x"00",x"00",x"0A",x"07",x"0A",x"3C",x"10",x"FE",x"A4",x"08",x"00",x"00",x"00",x"00",x"00",x"01",x"5A",x"F4",x"A8",x"60",x"00",x"00",x"00",x"FF",x"2D",x"1E",x"34",x"00",x"00",x"00",x"00",x"00",x"D2",x"E1",x"CB",x"FE",x"34",x"E2",x"40",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"18",x"3C",x"0E",x"03",x"06",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"B3",x"39",x"39",x"39",x"9B",x"C7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E7",x"C7",x"E7",x"E7",x"E7",x"E7",x"81",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"83",x"39",x"F1",x"C3",x"87",x"1F",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81",x"F3",x"E7",x"C3",x"F9",x"39",x"83",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E3",x"C3",x"93",x"33",x"01",x"F3",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"3F",x"03",x"F9",x"F9",x"39",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"9F",x"3F",x"03",x"39",x"39",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"39",x"F3",x"E7",x"CF",x"CF",x"CF",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"83",x"39",x"39",x"83",x"39",x"39",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"83",x"39",x"39",x"81",x"F9",x"F3",x"87",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"93",x"39",x"39",x"01",x"39",x"39",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"4A",x"2C",x"3E",x"78",x"3C",x"56",x"81",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"99",x"3F",x"3F",x"3F",x"99",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"33",x"39",x"39",x"39",x"33",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"3F",x"3F",x"03",x"3F",x"3F",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"3F",x"3F",x"03",x"3F",x"3F",x"3F",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C1",x"9F",x"3F",x"31",x"39",x"99",x"C1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"39",x"39",x"01",x"39",x"39",x"39",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81",x"E7",x"E7",x"E7",x"E7",x"E7",x"81",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"CF",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"83",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"81",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"11",x"01",x"01",x"29",x"39",x"39",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"19",x"09",x"01",x"21",x"31",x"39",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"83",x"39",x"39",x"39",x"39",x"39",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"39",x"39",x"39",x"03",x"3F",x"3F",x"FF",x"00",x"00",x"00",x"00",x"00",x"38",x"FF",x"FF",x"1F",x"3F",x"7F",x"7C",x"7C",x"00",x"44",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"39",x"39",x"31",x"07",x"23",x"31",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"33",x"3F",x"83",x"F9",x"39",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"39",x"39",x"39",x"39",x"39",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"39",x"39",x"11",x"83",x"C7",x"EF",x"FF",
																	x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"99",x"99",x"99",x"C3",x"E7",x"E7",x"E7",x"FF",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"FF",x"FF",x"EF",x"EF",x"EF",x"EF",x"EF",x"E7",x"00",x"FF",x"6F",x"2F",x"2F",x"2F",x"2F",x"2F",x"FD",x"FB",x"FB",x"F7",x"74",x"2F",x"8F",x"DF",x"02",x"06",x"04",x"0C",x"8F",x"D9",x"F0",x"70",x"DF",x"BF",x"BF",x"7F",x"F7",x"FA",x"F8",x"FC",x"20",x"60",x"40",x"C0",x"98",x"0D",x"0F",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",
																	x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"81",x"BD",x"A5",x"AD",x"A1",x"BF",x"80",x"FF",x"7E",x"42",x"5A",x"52",x"5E",x"40",x"7F",x"00",x"81",x"BD",x"A5",x"B5",x"85",x"FD",x"01",x"FF",x"7E",x"42",x"5A",x"4A",x"7A",x"02",x"FE",x"00",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",
																	x"00",x"00",x"00",x"00",x"07",x"07",x"0F",x"0F",x"00",x"00",x"00",x"00",x"07",x"07",x"0D",x"08",x"07",x"0F",x"07",x"67",x"C3",x"E4",x"CE",x"DE",x"02",x"00",x"00",x"00",x"02",x"07",x"09",x"11",x"FE",x"FE",x"7F",x"63",x"01",x"00",x"01",x"03",x"19",x"09",x"0C",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"3F",x"7F",x"7F",x"7C",x"78",x"F8",x"F8",
																	x"00",x"00",x"00",x"18",x"3C",x"3C",x"FF",x"FF",x"FC",x"FC",x"78",x"20",x"04",x"0C",x"78",x"F0",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"00",x"70",x"F8",x"F8",x"A0",x"20",x"20",x"40",x"F0",x"F8",x"FC",x"FC",x"F8",x"F8",x"F8",x"F0",x"F0",x"E0",x"E0",x"3C",x"CC",x"84",x"84",x"0C",x"0C",x"1C",x"FC",x"FC",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"FC",x"FC",x"F8",x"F8",x"F0",x"F0",x"F8",x"00",x"00",x"04",x"0E",x"0F",x"0F",x"FF",x"FF",x"7C",x"7C",x"38",x"30",x"01",x"03",x"1E",x"3C",x"07",x"07",x"0F",x"0F",x"07",x"0F",x"07",x"07",x"07",x"07",x"0D",x"08",x"02",x"00",x"00",x"00",x"01",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"07",x"07",x"07",x"07",
																	x"00",x"00",x"00",x"01",x"09",x"1F",x"1F",x"0F",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"03",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"0F",x"07",x"07",x"03",x"01",x"00",x"03",x"07",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"E0",x"E0",x"E0",x"A0",x"20",x"20",x"40",
																	x"C0",x"00",x"60",x"F0",x"F0",x"F8",x"F8",x"F8",x"40",x"E0",x"F0",x"F8",x"F8",x"F8",x"F8",x"C8",x"F8",x"70",x"70",x"F8",x"E0",x"E0",x"C0",x"00",x"88",x"88",x"88",x"08",x"18",x"18",x"38",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E0",x"E0",x"C0",x"80",x"80",x"80",x"C0",x"00",x"10",x"10",x"30",x"F0",x"E0",x"FF",x"FF",x"E0",x"F0",x"F0",x"D0",x"30",x"20",x"E0",x"C0",
																	x"00",x"0F",x"0F",x"1F",x"1F",x"0F",x"1F",x"0F",x"00",x"0F",x"0F",x"1B",x"11",x"05",x"00",x"00",x"0F",x"03",x"03",x"07",x"04",x"00",x"08",x"08",x"00",x"00",x"01",x"07",x"07",x"07",x"0F",x"0F",x"18",x"18",x"1C",x"1C",x"1C",x"F9",x"F2",x"E5",x"1F",x"1F",x"07",x"03",x"01",x"01",x"03",x"07",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"07",x"0F",x"0F",x"1F",x"1E",x"1E",x"3E",
																	x"00",x"00",x"08",x"1C",x"FC",x"7C",x"FF",x"FF",x"3E",x"1E",x"06",x"00",x"E0",x"7C",x"3C",x"08",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"80",x"C0",x"C0",x"C0",x"40",x"40",x"40",x"80",x"80",x"00",x"38",x"7C",x"7C",x"7E",x"7E",x"80",x"C0",x"F0",x"F8",x"FC",x"FC",x"FE",x"F8",x"3F",x"1F",x"07",x"03",x"7B",x"87",x"0E",x"0E",x"F0",x"F0",x"F8",x"F8",x"F8",x"F8",x"F0",x"F0",
																	x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"F8",x"F0",x"B0",x"78",x"F8",x"F8",x"7C",x"FF",x"FF",x"FF",x"9F",x"67",x"F2",x"F8",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"9F",x"0F",x"07",x"18",x"38",x"7C",x"F8",x"E0",x"C0",x"00",x"00",x"18",x"33",x"63",x"C7",x"E7",x"CF",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"F0",x"F8",x"FE",x"FF",x"FF",
																	x"00",x"00",x"00",x"07",x"07",x"06",x"00",x"00",x"3F",x"0F",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"06",x"0E",x"18",x"1B",x"3B",x"0B",x"00",x"03",x"07",x"0F",x"1F",x"0C",x"84",x"FC",x"09",x"04",x"0E",x"15",x"15",x"24",x"02",x"00",x"FE",x"FF",x"FF",x"7F",x"1F",x"3F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"1E",x"1E",x"1E",x"3E",x"3C",
																	x"00",x"00",x"00",x"00",x"00",x"18",x"FF",x"FF",x"3C",x"3C",x"7C",x"7C",x"38",x"00",x"22",x"3F",x"7C",x"7E",x"FE",x"FE",x"7E",x"FE",x"7E",x"7C",x"7C",x"7E",x"DE",x"8E",x"2A",x"02",x"02",x"04",x"5C",x"7C",x"7C",x"70",x"06",x"8F",x"9F",x"9F",x"40",x"C6",x"CE",x"FF",x"FF",x"7F",x"7F",x"6F",x"DF",x"FE",x"7C",x"38",x"10",x"80",x"00",x"00",x"27",x"02",x"80",x"C0",x"C0",x"80",x"80",x"80",
																	x"00",x"70",x"FF",x"DF",x"67",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"1F",x"1F",x"0F",x"1F",x"00",x"00",x"0F",x"0F",x"1B",x"11",x"05",x"00",x"0F",x"0F",x"FC",x"FE",x"FF",x"FF",x"7F",x"1E",x"00",x"00",x"3F",x"3F",x"7F",x"7F",x"7F",x"1F",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"07",x"07",x"07",x"03",x"03",x"03",x"03",
																	x"00",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"40",x"40",x"C0",x"80",x"00",x"10",x"18",x"0C",x"0C",x"0E",x"40",x"80",x"C0",x"F0",x"F8",x"FC",x"FC",x"FE",x"FE",x"FE",x"7F",x"63",x"01",x"00",x"00",x"00",x"19",x"09",x"0C",x"1C",x"3E",x"7F",x"FF",x"FB",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"E3",x"FC",x"FD",x"FB",x"7F",x"7F",x"3F",x"3F",x"1C",
																	x"00",x"00",x"00",x"0C",x"3E",x"78",x"FF",x"FF",x"01",x"03",x"07",x"03",x"21",x"61",x"F8",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"1F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FE",x"F8",x"E0",x"C0",x"00",x"00",x"0F",x"0F",x"03",x"1B",x"39",x"70",x"70",x"F0",x"00",x"00",x"00",x"1E",x"3F",x"7F",x"7F",x"FF",
																	x"F8",x"F0",x"F0",x"E4",x"FE",x"7F",x"0E",x"00",x"9F",x"07",x"07",x"1B",x"01",x"81",x"F1",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"80",x"C0",x"9C",x"3E",x"3E",x"3E",x"1E",x"40",x"80",x"78",x"FC",x"FE",x"FE",x"FE",x"FE",x"1F",x"1F",x"0F",x"0F",x"17",x"FE",x"7E",x"7C",x"F1",x"E0",x"F0",x"F0",x"F0",x"F0",x"81",x"83",
																	x"01",x"03",x"07",x"03",x"01",x"01",x"00",x"00",x"01",x"03",x"07",x"3E",x"7E",x"7E",x"FF",x"FF",x"01",x"02",x"02",x"02",x"00",x"00",x"00",x"08",x"F7",x"F7",x"FB",x"FB",x"F8",x"78",x"78",x"70",x"3C",x"3C",x"78",x"F0",x"00",x"00",x"00",x"00",x"04",x"0C",x"78",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"7E",x"FE",x"FE",x"00",x"00",x"00",x"00",x"7C",x"7E",x"DE",x"8E",
																	x"7E",x"FE",x"7E",x"7C",x"38",x"3C",x"78",x"00",x"2A",x"02",x"02",x"04",x"00",x"0C",x"7E",x"FF",x"07",x"07",x"0F",x"8F",x"8F",x"EF",x"EF",x"FF",x"FF",x"FF",x"FF",x"7F",x"7B",x"11",x"10",x"80",x"7E",x"5E",x"4C",x"40",x"00",x"00",x"00",x"00",x"80",x"E0",x"F0",x"FC",x"F8",x"F8",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F8",x"FC",x"7C",x"7C",x"7E",
																	x"00",x"02",x"07",x"07",x"03",x"03",x"02",x"02",x"3E",x"3C",x"19",x"09",x"01",x"03",x"02",x"02",x"00",x"00",x"00",x"01",x"01",x"03",x"07",x"03",x"00",x"00",x"00",x"01",x"01",x"03",x"07",x"3E",x"01",x"01",x"00",x"00",x"01",x"02",x"02",x"02",x"7E",x"7E",x"FF",x"FF",x"F7",x"F7",x"FB",x"FB",x"00",x"00",x"00",x"08",x"3C",x"3C",x"78",x"F0",x"F8",x"78",x"78",x"70",x"04",x"0C",x"78",x"F0",
																	x"80",x"C0",x"C0",x"E0",x"E0",x"E0",x"F0",x"60",x"80",x"80",x"80",x"80",x"98",x"DF",x"CF",x"5F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"0F",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"03",x"05",x"00",x"00",x"00",x"01",x"01",x"03",x"F3",x"FA",x"01",x"01",x"00",x"00",x"01",x"32",x"1A",x"1A",x"FE",x"FE",x"FF",x"7F",x"1F",x"0F",x"07",x"07",
																	x"38",x"3C",x"78",x"00",x"07",x"07",x"0F",x"8F",x"00",x"0C",x"7E",x"FF",x"FF",x"FF",x"FF",x"7F",x"8F",x"EF",x"EF",x"FF",x"7E",x"5E",x"4C",x"40",x"7B",x"11",x"10",x"80",x"80",x"E0",x"F0",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F8",x"F8",x"F0",x"F0",x"F0",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"02",x"07",x"07",x"FC",x"7C",x"7C",x"7E",x"3E",x"3C",x"19",x"09",
																	x"03",x"03",x"02",x"02",x"00",x"00",x"00",x"00",x"01",x"03",x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"7C",x"7E",x"FE",x"00",x"00",x"00",x"00",x"38",x"7C",x"7E",x"C4",x"FE",x"FF",x"3F",x"27",x"0F",x"02",x"00",x"00",x"94",x"A0",x"01",x"01",x"03",x"03",x"07",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"E0",x"E0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"E0",x"E0",x"B0",x"10",x"E0",x"F0",x"E0",x"E6",x"C3",x"27",x"73",x"7B",x"40",x"00",x"00",x"00",x"40",x"E0",x"90",x"88",x"7F",x"7F",x"FE",x"C6",x"80",x"00",x"80",x"C0",x"98",x"90",x"30",x"00",x"00",x"00",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"FC",x"FE",x"FE",x"3E",x"1E",x"1F",x"1F",
																	x"00",x"00",x"00",x"18",x"3C",x"3C",x"FF",x"FF",x"3F",x"3F",x"1E",x"04",x"20",x"30",x"1E",x"0F",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"07",x"07",x"07",x"07",x"03",x"00",x"0E",x"1F",x"1F",x"05",x"04",x"04",x"02",x"0F",x"1F",x"3F",x"3F",x"1F",x"1F",x"1F",x"0F",x"0F",x"07",x"07",x"3C",x"33",x"21",x"21",x"30",x"30",x"38",x"3F",x"3F",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"3F",x"3F",x"1F",x"1F",x"0F",x"0F",x"1F",x"00",x"00",x"20",x"70",x"F0",x"F0",x"FF",x"FF",x"3E",x"3E",x"1C",x"0C",x"80",x"C0",x"78",x"3C",x"E0",x"E0",x"F0",x"F0",x"E0",x"F0",x"E0",x"E0",x"E0",x"E0",x"B0",x"10",x"40",x"00",x"00",x"00",x"80",x"80",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",
																	x"00",x"00",x"00",x"80",x"90",x"F8",x"F8",x"F0",x"E0",x"C0",x"C0",x"80",x"00",x"00",x"00",x"C0",x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"C0",x"C0",x"E0",x"E0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"F0",x"E0",x"E0",x"C0",x"80",x"00",x"C0",x"E0",x"03",x"07",x"07",x"07",x"07",x"07",x"07",x"03",x"03",x"07",x"07",x"07",x"05",x"04",x"04",x"02",
																	x"03",x"00",x"06",x"0F",x"0F",x"1F",x"1F",x"1F",x"02",x"07",x"0F",x"1F",x"1F",x"1F",x"1F",x"13",x"1F",x"0E",x"0E",x"1F",x"07",x"07",x"03",x"00",x"11",x"11",x"11",x"10",x"18",x"18",x"1C",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"07",x"07",x"03",x"01",x"01",x"01",x"03",x"00",x"08",x"08",x"0C",x"0F",x"07",x"FF",x"FF",x"07",x"0F",x"0F",x"0B",x"0C",x"04",x"07",x"03",
																	x"00",x"F0",x"F0",x"F8",x"F8",x"F0",x"F8",x"F0",x"00",x"F0",x"F0",x"D8",x"88",x"A0",x"00",x"00",x"F0",x"C0",x"C0",x"E0",x"20",x"00",x"10",x"10",x"00",x"00",x"80",x"E0",x"E0",x"E0",x"F0",x"F0",x"18",x"18",x"38",x"38",x"38",x"9F",x"4F",x"A7",x"F8",x"F8",x"E0",x"C0",x"80",x"80",x"C0",x"E0",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"E0",x"F0",x"F0",x"F8",x"78",x"78",x"7C",
																	x"00",x"00",x"10",x"38",x"3F",x"3E",x"FF",x"FF",x"7C",x"78",x"60",x"00",x"07",x"3E",x"3C",x"10",x"00",x"01",x"03",x"03",x"03",x"03",x"03",x"03",x"00",x"01",x"03",x"03",x"03",x"02",x"02",x"02",x"01",x"01",x"00",x"1C",x"3E",x"3E",x"7E",x"7E",x"01",x"03",x"0F",x"1F",x"3F",x"3F",x"7F",x"1F",x"FC",x"F8",x"E0",x"C0",x"DE",x"E1",x"70",x"70",x"0F",x"0F",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",
																	x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"1F",x"0F",x"0D",x"1E",x"1F",x"1F",x"3E",x"E3",x"E1",x"02",x"06",x"04",x"0C",x"F9",x"00",x"2F",x"3D",x"FE",x"FE",x"FC",x"FC",x"F9",x"00",x"18",x"1C",x"3E",x"1F",x"07",x"03",x"00",x"00",x"18",x"CC",x"C6",x"E3",x"E7",x"F3",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"0F",x"1F",x"7F",x"FF",x"FF",
																	x"00",x"00",x"00",x"E0",x"E0",x"60",x"00",x"00",x"FC",x"F0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"60",x"70",x"18",x"D8",x"DC",x"D0",x"00",x"C0",x"E0",x"F0",x"F8",x"30",x"21",x"3F",x"90",x"20",x"70",x"A8",x"A8",x"24",x"40",x"00",x"7F",x"FF",x"FF",x"FE",x"F8",x"FC",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"78",x"78",x"78",x"7C",x"3C",
																	x"00",x"00",x"00",x"00",x"00",x"18",x"FF",x"FF",x"3C",x"3C",x"3E",x"3E",x"1C",x"00",x"44",x"FC",x"3E",x"7E",x"7F",x"7F",x"7E",x"7F",x"7E",x"3E",x"3E",x"7E",x"7B",x"71",x"54",x"40",x"40",x"20",x"3A",x"3E",x"3E",x"0E",x"60",x"F1",x"F9",x"F9",x"02",x"63",x"73",x"FF",x"FF",x"FE",x"FE",x"F6",x"FB",x"7F",x"3E",x"1C",x"08",x"01",x"00",x"00",x"E4",x"40",x"01",x"03",x"03",x"01",x"01",x"01",
																	x"00",x"0E",x"FF",x"FB",x"E6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F8",x"F8",x"F0",x"F8",x"00",x"00",x"F0",x"F0",x"D8",x"88",x"A0",x"00",x"F0",x"F0",x"3F",x"7F",x"FF",x"FF",x"FE",x"78",x"00",x"00",x"FC",x"FC",x"FE",x"FE",x"FE",x"F8",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"E0",x"E0",x"E0",x"C0",x"C0",x"C0",x"C0",
																	x"00",x"00",x"01",x"03",x"03",x"03",x"03",x"03",x"00",x"00",x"01",x"03",x"03",x"03",x"02",x"02",x"03",x"01",x"00",x"08",x"18",x"30",x"30",x"70",x"02",x"01",x"03",x"0F",x"1F",x"3F",x"3F",x"7F",x"7F",x"7F",x"FE",x"C6",x"80",x"00",x"00",x"00",x"98",x"90",x"30",x"38",x"7C",x"FE",x"FF",x"DF",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"C7",x"3F",x"BF",x"DF",x"FE",x"FE",x"FC",x"FC",x"38",
																	x"00",x"00",x"00",x"30",x"7C",x"1E",x"FF",x"FF",x"80",x"C0",x"E0",x"C0",x"84",x"86",x"1F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F8",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"7F",x"1F",x"07",x"03",x"00",x"00",x"F0",x"F0",x"C0",x"D8",x"9C",x"0E",x"0E",x"0F",x"00",x"00",x"00",x"78",x"FC",x"FE",x"FE",x"FF",
																	x"1F",x"0F",x"0F",x"27",x"7F",x"FE",x"70",x"00",x"F9",x"E0",x"E0",x"D8",x"80",x"81",x"8F",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"0F",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01",x"03",x"39",x"7C",x"7C",x"7C",x"78",x"02",x"01",x"1E",x"3F",x"7F",x"7F",x"7F",x"7F",x"F8",x"F8",x"F0",x"F0",x"E8",x"7F",x"7E",x"3E",x"8F",x"07",x"0F",x"0F",x"0F",x"0F",x"81",x"C1",
																	x"80",x"C0",x"E0",x"C0",x"80",x"80",x"00",x"00",x"80",x"C0",x"E0",x"7C",x"7E",x"7E",x"FF",x"FF",x"80",x"40",x"40",x"40",x"00",x"00",x"00",x"10",x"EF",x"EF",x"DF",x"DF",x"1F",x"1E",x"1E",x"0E",x"3C",x"3C",x"1E",x"0F",x"00",x"00",x"00",x"00",x"20",x"30",x"1E",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"7E",x"7F",x"7F",x"00",x"00",x"00",x"00",x"3E",x"7E",x"7B",x"71",
																	x"7E",x"7F",x"7E",x"3E",x"1C",x"3C",x"1E",x"00",x"54",x"40",x"40",x"20",x"00",x"30",x"7E",x"FF",x"E0",x"E0",x"F0",x"F1",x"F1",x"F7",x"F7",x"FF",x"FF",x"FF",x"FF",x"FE",x"DE",x"88",x"08",x"01",x"7E",x"7A",x"32",x"02",x"00",x"00",x"00",x"00",x"01",x"07",x"0F",x"3F",x"1F",x"1F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"1F",x"3F",x"3E",x"3E",x"7E",
																	x"00",x"40",x"E0",x"E0",x"C0",x"C0",x"40",x"40",x"7C",x"3C",x"98",x"90",x"80",x"C0",x"40",x"40",x"00",x"00",x"00",x"80",x"80",x"C0",x"E0",x"C0",x"00",x"00",x"00",x"80",x"80",x"C0",x"E0",x"7C",x"80",x"80",x"00",x"00",x"80",x"40",x"40",x"40",x"7E",x"7E",x"FF",x"FF",x"EF",x"EF",x"DF",x"DF",x"00",x"00",x"00",x"10",x"3C",x"3C",x"1E",x"0F",x"1F",x"1E",x"1E",x"0E",x"20",x"30",x"1E",x"0F",
																	x"01",x"03",x"03",x"07",x"07",x"07",x"0F",x"06",x"01",x"01",x"01",x"01",x"19",x"FB",x"F3",x"FA",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"F0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"C0",x"A0",x"00",x"00",x"00",x"80",x"80",x"C0",x"CF",x"5F",x"80",x"80",x"00",x"00",x"80",x"4C",x"58",x"58",x"7F",x"7F",x"FF",x"FE",x"F8",x"F0",x"E0",x"E0",
																	x"1C",x"3C",x"1E",x"00",x"E0",x"E0",x"F0",x"F1",x"00",x"30",x"7E",x"FF",x"FF",x"FF",x"FF",x"FE",x"F1",x"F7",x"F7",x"FF",x"7E",x"7A",x"32",x"02",x"DE",x"88",x"08",x"01",x"01",x"07",x"0F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"40",x"E0",x"E0",x"3F",x"3E",x"3E",x"7E",x"7C",x"3C",x"98",x"90",
																	x"C0",x"C0",x"40",x"40",x"00",x"00",x"00",x"00",x"80",x"C0",x"40",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"3E",x"7E",x"7F",x"00",x"00",x"00",x"00",x"1C",x"3E",x"7E",x"23",x"7F",x"FF",x"FC",x"E4",x"F0",x"40",x"00",x"00",x"29",x"05",x"80",x"80",x"C0",x"C0",x"E0",x"F0",x"00",x"00",x"30",x"70",x"70",x"60",x"60",x"C0",x"E0",x"E0",x"D0",x"90",x"30",x"20",x"60",x"C0",
																	x"67",x"EF",x"E7",x"C7",x"C3",x"CC",x"DC",x"FE",x"02",x"00",x"00",x"00",x"C2",x"CF",x"13",x"11",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"03",x"03",x"02",x"02",x"00",x"00",x"FF",x"FF",x"01",x"03",x"02",x"02",x"00",x"00",x"00",x"00",x"C0",x"C0",x"40",x"40",x"00",x"00",x"FF",x"FF",x"80",x"C0",x"40",x"40",x"00",x"00",x"00",x"00",
																	x"08",x"18",x"1C",x"18",x"1C",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"04",x"0E",x"06",x"00",x"01",x"01",x"02",x"00",x"18",x"39",x"F9",x"F9",x"00",x"01",x"03",x"07",x"1F",x"3F",x"1F",x"0F",x"FF",x"FF",x"DF",x"8F",x"2B",x"83",x"83",x"E7",x"C3",x"83",x"A1",x"F1",x"F5",x"FD",x"FD",x"FB",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"70",x"10",x"7F",x"7F",x"3F",x"00",x"03",x"0F",x"13",x"01",x"06",x"06",x"06",x"03",x"03",x"06",x"04",x"00",x"00",x"00",x"38",x"60",x"80",x"FE",x"FC",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"60",x"20",x"00",x"00",x"00",x"1C",x"06",x"01",x"7F",x"3F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",
																	x"C0",x"E0",x"F0",x"E0",x"40",x"F0",x"C0",x"C0",x"C0",x"E0",x"70",x"20",x"C0",x"00",x"00",x"00",x"07",x"0F",x"1F",x"0F",x"1F",x"3F",x"0F",x"1F",x"07",x"0F",x"1F",x"0E",x"1A",x"3A",x"08",x"1C",x"00",x"10",x"78",x"38",x"3C",x"1C",x"EF",x"FF",x"00",x"90",x"98",x"C8",x"CC",x"CC",x"0C",x"18",x"00",x"08",x"1E",x"1C",x"3C",x"38",x"F7",x"FF",x"00",x"09",x"19",x"13",x"33",x"33",x"30",x"18",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"3C",x"1E",x"1E",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"7E",x"3F",x"3F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
																	x"00",x"00",x"7E",x"3F",x"3F",x"00",x"00",x"3E",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1E",x"00",x"00",x"7E",x"3F",x"3F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"7F",x"7F",x"55",x"55",x"55",x"55",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"77",x"67",x"41",x"7F",x"7F",x"7F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
																	x"00",x"00",x"7E",x"3F",x"3F",x"0C",x"08",x"7E",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"16",x"24",x"7E",x"3F",x"3F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"18",x"1C",x"7E",x"3F",x"00",x"14",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"14",x"34",x"36",x"67",x"67",x"43",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"1F",x"09",x"14",x"36",x"13",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1D",x"1A",x"3E",x"14",x"0D",x"1F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"C0",x"94",x"B6",x"E4",x"C8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"DC",x"AC",x"BE",x"94",x"D8",x"FC",x"F8",x"00",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DD",x"77",x"AA",x"55",x"22",x"88",x"00",x"11",x"00",x"77",x"AA",x"55",x"22",x"88",x"00",x"11",x"00",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"EE",x"00",x"FF",x"FC",x"F5",x"F5",x"F5",x"F5",x"F5",x"CE",x"87",x"00",x"00",x"00",x"20",x"1F",x"00",x"F1",x"B8",x"7F",x"7F",x"3F",x"3F",x"1F",x"00",
																	x"00",x"00",x"00",x"08",x"04",x"06",x"03",x"00",x"0F",x"07",x"07",x"1F",x"3F",x"7F",x"FF",x"FB",x"00",x"00",x"00",x"10",x"20",x"60",x"C0",x"00",x"F0",x"E0",x"E0",x"F8",x"FC",x"FE",x"FF",x"DF",x"78",x"30",x"00",x"00",x"0C",x"0C",x"FF",x"FF",x"07",x"0F",x"1F",x"3E",x"32",x"10",x"26",x"3F",x"1E",x"0C",x"00",x"00",x"30",x"30",x"FF",x"FF",x"E0",x"F0",x"F8",x"7C",x"4C",x"08",x"64",x"FC",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"11",x"83",x"C7",x"83",x"11",x"39",x"FF",x"FF",x"FC",x"E0",x"60",x"30",x"18",x"FF",x"FF",x"FF",x"FC",x"D8",x"7C",x"3E",x"1F",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"39",x"39",x"03",x"39",x"39",x"03",x"FF",x"FF",x"FF",x"03",x"06",x"0C",x"18",x"FF",x"FF",x"FF",x"FF",x"1F",x"3E",x"7C",x"F8",x"00",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"60",x"F0",x"F0",x"F8",x"F8",x"F8",x"40",x"E0",x"F0",x"F8",x"F8",x"FC",x"FC",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF");
																		
	
	constant DUCK_HUNT_CHR_ROM : CHR_ROM_ARRAY := (x"00",x"00",x"00",x"01",x"02",x"03",x"03",x"05",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"60",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"20",x"60",x"E0",x"60",x"E0",x"E0",x"E0",x"00",x"00",x"00",x"04",x"0E",x"0E",x"0E",x"0E",x"00",x"00",x"00",x"1A",x"31",x"71",x"75",x"75",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"E0",x"E0",x"C0",x"80",
																	x"07",x"07",x"07",x"03",x"03",x"01",x"01",x"00",x"03",x"03",x"03",x"01",x"01",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F9",x"FB",x"F7",x"CF",x"BF",x"F0",x"F0",x"F0",x"F8",x"FB",x"FF",x"FF",x"FF",x"04",x"00",x"00",x"C1",x"E3",x"EF",x"DF",x"FE",x"7B",x"7F",x"FE",x"3D",x"93",x"CE",x"DC",x"F8",x"1E",x"7C",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"1E",x"60",x"C0",x"80",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"01",x"01",x"01",x"03",x"0F",x"00",x"00",x"00",x"01",x"01",x"01",x"03",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"F8",x"FC",x"FC",x"F8",x"F0",x"E0",x"C0",x"00",x"00",x"F8",x"F0",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"06",x"0E",x"0E",x"04",x"00",x"00",
																	x"FE",x"FC",x"F0",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"08",x"38",x"70",x"F0",x"F0",x"60",x"00",x"00",x"04",x"0E",x"0E",x"0E",x"0E",x"04",x"00",x"00",x"1A",x"31",x"71",x"75",x"75",x"7B",x"00",x"50",x"70",x"38",x"3C",x"7C",x"78",x"F8",x"00",x"50",x"70",x"30",x"21",x"63",x"67",x"E7",x"00",x"00",x"00",x"1F",x"FF",x"7F",x"0F",x"07",x"00",x"00",x"00",x"1F",x"3F",x"07",x"03",x"03",
																	x"00",x"00",x"01",x"03",x"C7",x"EF",x"DF",x"BF",x"00",x"00",x"00",x"03",x"C7",x"FF",x"FF",x"FF",x"00",x"00",x"C0",x"E0",x"E0",x"C0",x"E0",x"FF",x"7F",x"FE",x"3C",x"90",x"C0",x"C0",x"E0",x"FF",x"03",x"03",x"01",x"01",x"01",x"03",x"0F",x"07",x"01",x"01",x"01",x"01",x"01",x"03",x"0F",x"02",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"E0",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"C7",x"03",x"00",x"FF",x"FF",x"FF",x"FF",x"C7",x"01",x"00",x"00",x"C0",x"F0",x"F8",x"FC",x"FF",x"EE",x"B0",x"C0",x"C0",x"F0",x"F8",x"FC",x"EE",x"A0",x"00",x"00",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"0E",x"0E",x"04",x"00",x"00",x"00",x"FC",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"38",x"70",x"F0",x"F0",x"60",x"00",
																	x"00",x"04",x"0E",x"0E",x"0E",x"0E",x"04",x"00",x"00",x"1A",x"31",x"71",x"75",x"75",x"7B",x"7F",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"67",x"B3",x"B0",x"D0",x"F0",x"F8",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"00",x"01",x"03",x"07",x"0F",x"BF",x"7F",x"FF",x"00",x"00",x"03",x"07",x"3F",x"FF",x"FF",x"FF",
																	x"00",x"C0",x"E0",x"E0",x"C0",x"C0",x"80",x"80",x"FE",x"3C",x"90",x"C0",x"C0",x"C0",x"80",x"80",x"07",x"07",x"0D",x"1D",x"33",x"0F",x"07",x"03",x"06",x"05",x"09",x"11",x"03",x"0F",x"02",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F3",x"E5",x"01",x"C0",x"C0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"C0",x"C0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",
																	x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"0E",x"0E",x"04",x"00",x"00",x"00",x"00",x"F3",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"09",x"38",x"70",x"F0",x"F0",x"60",x"00",x"00",x"F0",x"F8",x"F8",x"F8",x"FC",x"FC",x"7E",x"1E",x"F0",x"F8",x"F8",x"78",x"7C",x"3C",x"0E",x"02",x"18",x"38",x"3C",x"3C",x"3E",x"5E",x"7F",x"7F",x"18",x"18",x"1C",x"1C",x"1E",x"0E",x"3F",x"3F",
																	x"3F",x"3F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"1F",x"1F",x"0F",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"01",x"03",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"00",x"00",x"03",x"03",x"83",x"C3",x"E7",x"FF",x"0F",x"0F",x"04",x"01",x"83",x"C3",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"2F",x"1F",x"1F",x"FF",x"FF",x"FF",x"FF",x"3F",x"0F",x"1F",x"1F",
																	x"1F",x"1F",x"1F",x"0F",x"07",x"03",x"00",x"00",x"1F",x"0E",x"04",x"00",x"08",x"1C",x"1C",x"0C",x"00",x"0F",x"3F",x"FF",x"FF",x"BF",x"7F",x"19",x"00",x"0F",x"3F",x"FF",x"7F",x"3F",x"19",x"00",x"00",x"01",x"03",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"0F",x"00",x"03",x"03",x"03",x"03",x"83",x"E7",x"FF",x"0F",x"04",x"01",x"03",x"03",x"83",x"E7",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"6F",x"1F",x"1F",x"1F",x"FF",x"FF",x"FF",x"7F",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"07",x"03",x"00",x"00",x"00",x"0E",x"04",x"00",x"08",x"1C",x"1C",x"1C",x"0C",x"00",x"00",x"01",x"01",x"03",x"07",x"0F",x"00",x"00",x"00",x"01",x"01",x"03",x"06",x"08",x"00",x"01",x"03",x"04",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"03",x"07",x"0F",x"0F",x"0F",x"0E",
																	x"03",x"03",x"03",x"03",x"03",x"07",x"0F",x"1F",x"04",x"01",x"03",x"03",x"03",x"07",x"0F",x"1F",x"3F",x"3F",x"77",x"6F",x"FF",x"FF",x"FF",x"FF",x"3F",x"3F",x"7F",x"7F",x"FF",x"DF",x"DF",x"8E",x"DF",x"8F",x"07",x"03",x"00",x"00",x"00",x"00",x"04",x"00",x"08",x"1C",x"1C",x"1C",x"0C",x"00",x"00",x"40",x"60",x"30",x"00",x"00",x"00",x"01",x"00",x"40",x"60",x"30",x"00",x"00",x"00",x"01",
																	x"80",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"80",x"00",x"00",x"00",x"00",x"00",x"C0",x"F1",x"0C",x"1E",x"1F",x"3F",x"3F",x"3F",x"3E",x"1E",x"00",x"00",x"00",x"00",x"0C",x"4C",x"C1",x"E1",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"3C",x"7C",x"F8",x"E0",x"03",x"07",x"0F",x"0F",x"1F",x"1F",x"1D",x"18",x"03",x"07",x"0F",x"0F",x"1D",x"1C",x"10",x"00",
																	x"F8",x"FC",x"FC",x"FC",x"FE",x"BE",x"1E",x"0F",x"F9",x"FD",x"FD",x"BC",x"3E",x"1E",x"0E",x"07",x"0C",x"00",x"00",x"00",x"00",x"40",x"F8",x"F0",x"F3",x"FF",x"FF",x"FF",x"7E",x"3C",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"E0",x"70",x"10",x"00",x"00",x"00",x"07",x"07",x"43",x"C3",x"87",x"07",x"07",x"07",x"03",x"03",x"43",x"C3",x"87",x"06",x"04",x"04",
																	x"FB",x"FF",x"FF",x"FF",x"FF",x"FC",x"FC",x"FC",x"FB",x"FF",x"FF",x"C7",x"04",x"00",x"00",x"00",x"E1",x"F3",x"F8",x"FC",x"FC",x"7C",x"1C",x"18",x"E1",x"F3",x"F8",x"FC",x"7C",x"1C",x"08",x"00",x"1F",x"03",x"07",x"07",x"06",x"00",x"00",x"00",x"F0",x"EC",x"F8",x"70",x"36",x"00",x"00",x"00",x"E0",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"06",x"6F",x"3E",x"1C",x"18",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"00",x"03",x"17",x"3F",x"7F",x"FE",x"FE",x"FC",x"00",x"03",x"17",x"3B",x"53",x"86",x"06",x"04",x"03",x"03",x"03",x"07",x"07",x"07",x"07",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"FC",x"F8",x"F8",x"F8",x"F8",x"F0",x"F3",x"FF",x"0C",x"08",x"08",x"08",x"18",x"10",x"12",x"1E",
																	x"00",x"00",x"04",x"0E",x"0E",x"0E",x"0E",x"04",x"00",x"00",x"1A",x"31",x"73",x"F3",x"F1",x"FB",x"00",x"17",x"0F",x"07",x"03",x"01",x"01",x"00",x"00",x"17",x"0F",x"03",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"F8",x"F8",x"F8",x"F8",x"70",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FC",x"F8",x"F0",x"C0",x"3E",x"3E",x"3F",x"0F",x"00",x"00",x"00",x"00",
																	x"00",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"FF",x"7E",x"40",x"00",x"00",x"00",x"00",x"00",x"7F",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"F8",x"F0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"F0",x"F8",x"F8",x"00",x"00",x"00",x"00",x"80",x"00",x"18",x"20",x"22",x"24",x"3C",x"00",x"E0",x"F0",x"F8",x"F8",x"FE",x"FC",x"F8",
																	x"7C",x"3D",x"3B",x"27",x"2F",x"1F",x"1F",x"1F",x"C8",x"C4",x"DC",x"F9",x"F0",x"E4",x"E0",x"E0",x"3F",x"3F",x"3F",x"3F",x"3C",x"00",x"FF",x"F8",x"CC",x"CA",x"C8",x"C0",x"40",x"00",x"FF",x"F8",x"00",x"00",x"00",x"00",x"00",x"30",x"78",x"78",x"00",x"00",x"00",x"00",x"00",x"30",x"68",x"70",x"F8",x"F0",x"F8",x"F8",x"F8",x"F8",x"F8",x"F0",x"78",x"70",x"30",x"00",x"00",x"90",x"00",x"00",
																	x"F0",x"E0",x"C0",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"80",x"40",x"30",x"08",x"04",x"04",x"E0",x"F0",x"78",x"3C",x"0E",x"07",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"07",x"07",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60",x"70",x"FE",x"FF",x"FF",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"00",x"E0",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",
																	x"00",x"07",x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"00",x"07",x"0F",x"0F",x"1F",x"3F",x"FF",x"FF",x"00",x"80",x"00",x"18",x"20",x"20",x"22",x"3C",x"00",x"E0",x"F0",x"F8",x"F8",x"F8",x"FE",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"1F",x"3F",x"7F",x"7F",x"7F",x"7C",x"78",x"01",x"02",x"04",x"0F",x"3F",x"1F",x"1F",x"0F",x"FE",x"FD",x"FB",x"F0",x"C0",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"80",x"C0",x"64",x"34",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1B",x"0B",x"04",x"04",x"04",x"04",x"04",x"04",x"06",x"06",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"3E",x"3E",x"3E",x"7E",x"7E",x"7E",x"7E",x"7E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7C",x"3C",x"3D",x"13",x"2F",x"0F",x"1F",x"1F",x"C8",x"C0",x"CE",x"FC",x"F0",x"F0",x"E2",x"E0",
																	x"0C",x"1E",x"FE",x"FE",x"FC",x"FC",x"FC",x"FC",x"0C",x"1A",x"3C",x"3E",x"9C",x"00",x"40",x"10",x"00",x"00",x"00",x"00",x"20",x"C0",x"00",x"FF",x"78",x"78",x"F8",x"F8",x"F8",x"F0",x"E0",x"FF",x"0E",x"0F",x"0F",x"0F",x"07",x"07",x"3F",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"FF",x"1E",x"06",x"87",x"E7",x"F7",x"F7",x"F1",x"FF",x"01",x"01",x"00",x"00",x"40",x"20",x"21",x"FF",
																	x"02",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"FE",x"FF",x"FC",x"FE",x"7F",x"3F",x"1F",x"9F",x"FF",x"7E",x"7E",x"3E",x"06",x"00",x"10",x"08",x"08",x"FF",x"7F",x"3F",x"FE",x"FC",x"FE",x"FE",x"FE",x"3F",x"3F",x"3F",x"3F",x"3F",x"3C",x"FF",x"FC",x"C1",x"C0",x"CC",x"CE",x"4C",x"00",x"FF",x"FC",x"F8",x"F8",x"F0",x"E0",x"00",x"00",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"0C",x"06",x"06",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"0E",x"1E",x"3C",x"78",x"70",x"70",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"0F",x"0F",x"0F",x"07",x"03",x"00",x"02",x"0C",x"3E",x"3B",x"01",x"00",x"00",x"00",x"FD",x"F3",x"C1",x"C0",x"E0",x"F0",x"F0",x"F8",x"00",x"00",x"00",x"00",x"80",x"C4",x"64",x"34",x"FF",x"FF",x"FF",x"FF",x"7F",x"3B",x"1B",x"0B",x"04",x"04",x"04",x"04",x"04",x"04",x"02",x"0A",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",
																	x"01",x"01",x"01",x"00",x"00",x"00",x"01",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"00",x"90",x"90",x"A6",x"CF",x"7F",x"FF",x"FF",x"F8",x"78",x"78",x"78",x"34",x"02",x"82",x"FF",x"1C",x"06",x"02",x"02",x"02",x"00",x"0F",x"FF",x"03",x"01",x"01",x"01",x"01",x"01",x"0F",x"FF",x"0A",x"0F",x"07",x"00",x"00",x"00",x"00",x"F0",x"F7",x"F0",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"7E",x"FE",x"FE",x"3E",x"1C",x"40",x"2F",x"2F",x"FF",x"7F",x"3F",x"FE",x"FC",x"F0",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"07",x"07",x"07",x"03",x"03",x"03",x"03",x"02",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"80",x"81",x"81",x"81",x"00",x"00",x"FF",x"FF",x"7F",x"7E",x"7E",x"7C",x"7C",x"3E",x"40",x"40",x"80",x"02",x"02",x"C2",x"64",x"34",x"BF",x"BF",x"7F",x"FD",x"FD",x"3D",x"1B",x"0B",x"04",x"04",x"04",x"04",x"04",x"04",x"12",x"12",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"0F",x"1F",x"1F",x"1F",x"1E",x"0C",x"00",x"0F",x"00",x"00",x"00",x"04",x"08",x"00",x"00",x"0F",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"FC",x"3E",x"1E",x"1F",x"0F",x"0F",x"07",x"3F",x"FF",x"1C",x"00",x"00",x"00",x"00",x"40",x"2E",x"2F",x"03",x"07",x"07",x"07",x"E7",x"F3",x"FF",x"FF",x"12",x"26",x"3F",x"0F",x"00",x"04",x"02",x"C2",x"EF",x"D8",x"C0",x"F0",x"FF",x"FF",x"FF",x"FF",x"7E",x"7E",x"3E",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"3E",x"1C",x"82",x"82",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"03",x"07",x"1F",x"1F",x"1F",x"1F",x"1F",x"01",x"01",x"02",x"03",x"01",x"18",x"7E",x"7F",x"FE",x"FE",x"FD",x"FC",x"F8",x"E0",x"80",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"62",x"32",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1D",x"0D",x"04",x"04",x"04",x"04",x"04",x"04",x"0A",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F2",
																	x"3E",x"3E",x"3E",x"7E",x"7E",x"7E",x"7E",x"1E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"0F",x"0F",x"0F",x"0F",x"07",x"07",x"03",x"0F",x"1F",x"0F",x"07",x"06",x"00",x"20",x"17",x"17",x"02",x"02",x"04",x"80",x"F0",x"F8",x"FF",x"FF",x"1E",x"06",x"00",x"00",x"00",x"00",x"03",x"FF",x"01",x"01",x"01",x"01",x"00",x"00",x"03",x"FF",
																	x"00",x"08",x"00",x"00",x"00",x"01",x"87",x"FF",x"F9",x"F7",x"FF",x"FF",x"FF",x"FE",x"F8",x"FE",x"0E",x"26",x"16",x"0E",x"3E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"DC",x"00",x"02",x"02",x"0F",x"1F",x"13",x"27",x"26",x"2E",x"4E",x"4C",x"0F",x"1F",x"1F",x"3B",x"3A",x"36",x"76",x"74",x"00",x"00",x"1E",x"3F",x"3F",x"7E",x"78",x"70",x"00",x"00",x"1E",x"3F",x"3F",x"7E",x"78",x"70",
																	x"4C",x"4C",x"4E",x"2E",x"1F",x"17",x"0B",x"07",x"74",x"74",x"76",x"36",x"13",x"18",x"0D",x"07",x"70",x"20",x"03",x"67",x"E7",x"CF",x"CF",x"8F",x"70",x"3E",x"3F",x"7C",x"FC",x"F8",x"F9",x"F9",x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"40",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"01",x"01",x"01",x"01",x"03",x"07",x"0F",x"3F",
																	x"0F",x"0F",x"0F",x"07",x"07",x"03",x"05",x"03",x"F8",x"F8",x"F8",x"FC",x"FD",x"FE",x"FE",x"FC",x"C0",x"C1",x"CF",x"BF",x"7F",x"FF",x"FF",x"FF",x"80",x"01",x"41",x"C0",x"88",x"02",x"10",x"00",x"F0",x"F8",x"F8",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"C8",x"E8",x"F0",x"00",x"00",x"00",x"80",x"04",x"04",x"04",x"06",x"02",x"02",x"03",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"07",x"0F",x"0F",x"1F",x"1F",x"1F",x"0F",x"4F",x"F8",x"F0",x"F3",x"E3",x"E3",x"E3",x"F3",x"C1",x"FF",x"FF",x"FF",x"EF",x"C0",x"80",x"80",x"80",x"04",x"00",x"00",x"E0",x"C0",x"80",x"80",x"80",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"09",x"0A",x"0C",x"08",x"00",x"00",x"00",x"FF",x"F6",x"F4",x"F0",x"F0",x"F8",x"F8",x"FC",
																	x"CE",x"87",x"07",x"03",x"00",x"00",x"00",x"00",x"C1",x"81",x"01",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F8",x"F8",x"F8",x"F8",x"70",x"00",x"40",x"20",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"FE",x"FC",x"FE",x"FE",x"7F",x"3F",x"1F",x"9F",x"FF",x"00",x"00",x"00",x"00",x"00",x"08",x"05",x"05",x"00",x"00",x"00",x"F8",x"FC",x"FE",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"F0",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"00",x"00",x"00",x"07",x"0F",x"1F",x"1F",x"FF",x"00",x"00",x"00",x"07",x"03",x"00",x"00",x"E0",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"F0",x"F8",x"F8",x"F8",x"70",x"00",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"F8",x"F0",x"E0",x"40",x"00",x"00",x"00",x"00",x"00",x"F0",x"F8",x"F8",x"F3",x"FF",x"FF",x"00",x"00",x"F0",x"F8",x"F8",x"D2",x"1E",x"1E",x"FF",x"FF",x"FF",x"FC",x"F8",x"F0",x"C0",x"00",x"3E",x"3F",x"3F",x"0C",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"0F",x"7F",x"FF",x"00",x"00",x"00",x"00",x"00",x"0F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"0F",x"FF",x"FF",x"FF",x"FF",x"37",x"07",x"03",x"13",x"03",x"03",x"03",x"01",x"01",x"00",x"00",x"00",x"FB",x"F1",x"E1",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E3",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"E2",x"FE",x"FE",x"FE",
																	x"FF",x"FF",x"FC",x"F8",x"F0",x"F0",x"F0",x"F8",x"FF",x"FF",x"FC",x"F0",x"F0",x"F0",x"F0",x"F8",x"F8",x"F8",x"F8",x"FC",x"FC",x"FC",x"3E",x"0E",x"F8",x"F8",x"F8",x"FC",x"BC",x"2C",x"0E",x"06",x"FE",x"FE",x"7E",x"7C",x"3C",x"38",x"38",x"38",x"F8",x"F8",x"7A",x"7C",x"3C",x"38",x"38",x"00",x"00",x"00",x"00",x"00",x"20",x"3A",x"3E",x"3F",x"00",x"00",x"00",x"00",x"20",x"30",x"38",x"3A",
																	x"3F",x"1F",x"1F",x"0F",x"0F",x"07",x"03",x"01",x"3F",x"1F",x"1F",x"0F",x"0F",x"07",x"03",x"01",x"00",x"03",x"07",x"05",x"01",x"0B",x"0F",x"0F",x"03",x"00",x"00",x"02",x"06",x"04",x"00",x"00",x"1E",x"1E",x"1E",x"3E",x"3C",x"18",x"00",x"00",x"01",x"01",x"01",x"05",x"0B",x"2E",x"18",x"00",x"20",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"10",x"18",x"38",x"38",x"38",x"1C",x"1C",x"1E",
																	x"11",x"10",x"08",x"04",x"02",x"01",x"00",x"00",x"0E",x"0F",x"07",x"0B",x"0D",x"1E",x"1F",x"1F",x"04",x"05",x"06",x"07",x"03",x"00",x"00",x"40",x"9B",x"DA",x"D9",x"F8",x"FC",x"FF",x"FF",x"BF",x"41",x"62",x"3C",x"00",x"00",x"00",x"00",x"00",x"BE",x"9C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"78",x"7C",x"00",x"00",x"00",x"00",x"00",x"30",x"78",x"7C",
																	x"7C",x"1C",x"0E",x"0E",x"06",x"04",x"00",x"00",x"7C",x"1C",x"0E",x"0E",x"07",x"07",x"03",x"07",x"00",x"00",x"07",x"08",x"00",x"00",x"00",x"3C",x"07",x"07",x"07",x"0F",x"0F",x"1F",x"3F",x"43",x"03",x"80",x"00",x"00",x"00",x"00",x"00",x"03",x"FC",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"04",x"58",x"CB",x"FB",x"FA",x"FA",x"02",x"07",x"FB",x"A7",x"34",x"04",x"05",x"05",x"05",x"00",
																	x"07",x"07",x"07",x"0F",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"0D",x"05",x"03",x"00",x"00",x"38",x"3C",x"3A",x"18",x"1C",x"0C",x"00",x"00",x"38",x"34",x"36",x"16",x"1A",x"0B",x"0E",x"06",x"06",x"07",x"0F",x"1E",x"0C",x"00",x"0D",x"05",x"05",x"F4",x"FD",x"FE",x"FE",x"FE",x"01",x"00",x"E0",x"18",x"04",x"02",x"02",x"01",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",
																	x"00",x"80",x"00",x"00",x"10",x"1C",x"0E",x"1B",x"FE",x"7F",x"FF",x"FF",x"EF",x"E3",x"F1",x"E0",x"80",x"40",x"20",x"A0",x"A0",x"80",x"88",x"88",x"70",x"B8",x"D8",x"58",x"58",x"78",x"70",x"70",x"90",x"90",x"A0",x"80",x"80",x"00",x"00",x"00",x"60",x"60",x"40",x"40",x"C0",x"C0",x"80",x"00",x"80",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"80",x"80",x"40",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"80",x"80",x"10",x"18",x"20",x"C0",x"00",x"70",x"78",x"78",x"E8",x"E0",x"C0",x"00",x"00",x"00",x"1C",x"3E",x"7F",x"07",x"03",x"07",x"00",x"00",x"1C",x"3E",x"7F",x"07",x"03",x"F7",x"1C",x"3E",x"3E",x"0F",x"07",x"07",x"07",x"C6",x"1C",x"3E",x"3E",x"0F",x"07",x"07",x"FF",x"FE",x"00",x"00",x"00",x"00",x"0C",x"07",x"00",x"00",x"00",x"01",x"0F",x"0F",x"03",x"00",x"00",x"00",
																	x"00",x"01",x"00",x"3C",x"C3",x"00",x"00",x"00",x"39",x"FE",x"FF",x"C3",x"0C",x"1F",x"1F",x"1F",x"03",x"00",x"00",x"00",x"00",x"80",x"00",x"03",x"FC",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FC",x"32",x"CA",x"24",x"02",x"01",x"01",x"00",x"00",x"FE",x"3E",x"DE",x"FF",x"FF",x"FF",x"FF",x"FF",x"88",x"44",x"24",x"A4",x"A6",x"8B",x"89",x"88",x"77",x"BB",x"DB",x"5B",x"59",x"70",x"70",x"70",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"C0",x"80",x"80",x"80",x"C0",x"E0",x"E0",x"40",x"00",x"00",x"00",x"00",x"01",x"07",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"01",x"07",x"0F",x"1F",x"1F",x"3E",x"3E",x"3E",x"3C",x"1C",x"1C",x"0C",x"00",x"3E",x"3E",x"3E",x"3C",x"1C",x"1C",x"0C",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"10",x"03",x"07",x"0F",x"0F",x"1F",x"1F",x"1F",x"0F",
																	x"10",x"10",x"08",x"08",x"08",x"04",x"03",x"00",x"0F",x"0F",x"07",x"07",x"07",x"03",x"00",x"00",x"C0",x"F0",x"F6",x"2E",x"1E",x"1E",x"1E",x"1E",x"C6",x"FF",x"FF",x"39",x"31",x"35",x"33",x"31",x"0F",x"77",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3B",x"0F",x"02",x"49",x"00",x"04",x"91",x"42",x"FF",x"FF",x"7F",x"3F",x"9F",x"C7",x"70",x"1F",x"3C",x"44",x"EE",x"C4",x"E0",x"F8",x"FF",x"FF",
																	x"0E",x"01",x"00",x"01",x"00",x"E8",x"B5",x"9E",x"F1",x"FE",x"FF",x"FF",x"FF",x"1F",x"4E",x"63",x"80",x"80",x"C0",x"40",x"40",x"40",x"40",x"40",x"7F",x"7F",x"3F",x"3F",x"3F",x"3F",x"3F",x"3F",x"FF",x"FF",x"F3",x"C9",x"C1",x"A1",x"10",x"80",x"3C",x"22",x"7F",x"3F",x"3F",x"7F",x"FF",x"FF",x"60",x"18",x"84",x"82",x"83",x"81",x"01",x"01",x"9F",x"E7",x"7B",x"7D",x"FC",x"7E",x"FE",x"FE",
																	x"80",x"C6",x"FE",x"FE",x"FE",x"7C",x"18",x"00",x"80",x"C6",x"FE",x"FE",x"FE",x"7C",x"18",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"F8",x"F8",x"FC",x"C0",x"20",x"04",x"04",x"0C",x"08",x"98",x"70",x"FC",x"FC",x"F8",x"F8",x"F0",x"F0",x"60",x"00",x"00",x"C0",x"E0",x"F0",x"76",x"2E",x"1E",x"1E",x"00",x"C0",x"E6",x"FF",x"7F",x"39",x"31",x"35",
																	x"1E",x"1E",x"0F",x"77",x"FF",x"FF",x"FF",x"FF",x"33",x"31",x"3B",x"0F",x"02",x"49",x"00",x"04",x"FF",x"FF",x"FF",x"7F",x"3F",x"8F",x"60",x"1F",x"91",x"42",x"3C",x"C4",x"C4",x"F0",x"FF",x"FF",x"FF",x"FF",x"F3",x"C9",x"C1",x"A1",x"10",x"00",x"89",x"42",x"3E",x"7F",x"7F",x"7F",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"02",x"01",x"03",x"07",x"0F",x"1F",x"1E",x"3C",x"3C",
																	x"0E",x"00",x"02",x"0E",x"06",x"44",x"3C",x"00",x"70",x"7C",x"7C",x"78",x"7C",x"38",x"10",x"00",x"C0",x"F0",x"F6",x"2E",x"1E",x"1E",x"1E",x"1E",x"C6",x"FF",x"FF",x"39",x"31",x"33",x"33",x"31",x"0F",x"77",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"3B",x"0F",x"02",x"49",x"00",x"04",x"11",x"43",x"3F",x"1F",x"5F",x"4F",x"27",x"10",x"4F",x"C0",x"7F",x"7F",x"FD",x"F8",x"F8",x"FF",x"BF",x"3F",
																	x"C0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"3F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"FD",x"F9",x"FA",x"F2",x"E4",x"08",x"F1",x"03",x"FF",x"FF",x"3F",x"9F",x"1F",x"FF",x"FE",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"03",x"0F",x"1F",x"7F",x"FE",x"02",x"04",x"08",x"30",x"61",x"C1",x"81",x"83",x"FC",x"F8",x"F0",x"C0",x"81",x"01",x"01",x"03",
																	x"03",x"07",x"07",x"0D",x"00",x"00",x"00",x"00",x"03",x"06",x"04",x"08",x"00",x"00",x"00",x"00",x"0C",x"1E",x"1E",x"1E",x"0C",x"00",x"00",x"00",x"3C",x"7E",x"FF",x"E9",x"F3",x"7F",x"7E",x"38",x"08",x"08",x"48",x"30",x"28",x"00",x"24",x"7E",x"74",x"F6",x"BE",x"DE",x"DC",x"FC",x"FC",x"7E",x"7E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"F8",x"7E",x"FD",x"FC",x"FC",x"EC",x"D8",x"DB",x"B7",
																	x"F8",x"F8",x"7C",x"3C",x"38",x"70",x"50",x"00",x"37",x"77",x"63",x"21",x"30",x"70",x"50",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"F0",x"E0",x"80",x"C0",x"40",x"00",x"00",x"80",x"80",x"80",x"80",x"80",x"00",x"00",x"00",x"20",x"30",x"30",x"30",x"F0",x"20",x"00",x"00",x"07",x"3F",x"7F",x"FF",x"FF",x"7F",x"1F",x"03",x"00",x"00",x"00",x"00",x"80",x"60",x"1C",x"03",
																	x"00",x"00",x"07",x"1F",x"3F",x"3F",x"1F",x"07",x"00",x"00",x"00",x"00",x"00",x"20",x"18",x"07",x"00",x"00",x"00",x"00",x"04",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"00",x"7E",x"FF",x"FF",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"C3",x"3C",x"00",x"00",
																	x"00",x"00",x"38",x"7C",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"1F",x"3F",x"7F",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"FF",x"FF",x"FF",x"7F",x"1F",x"07",x"00",x"00",x"00",x"00",x"80",x"60",x"1C",x"07",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"C3",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"F8",x"E0",x"80",x"80",x"C0",x"60",x"00",x"00",x"07",x"04",x"04",x"07",x"01",x"05",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"07",x"05",x"05",x"02",x"05",x"05",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"27",x"25",x"25",x"25",x"25",x"25",x"27",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"27",x"24",x"24",x"27",x"21",x"25",x"27",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"27",x"24",x"24",x"27",x"25",x"25",x"27",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"77",x"55",x"15",x"35",x"65",x"45",x"77",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"75",x"55",x"15",x"37",x"61",x"41",x"71",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"77",x"15",x"15",x"75",x"15",x"15",x"77",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"77",x"55",x"55",x"55",x"55",x"55",x"77",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"C7",x"B3",x"39",x"39",x"39",x"9B",x"C7",x"FF",x"38",x"4C",x"C6",x"C6",x"C6",x"64",x"38",x"00",x"E7",x"C7",x"E7",x"E7",x"E7",x"E7",x"81",x"FF",x"18",x"38",x"18",x"18",x"18",x"18",x"7E",x"00",x"83",x"39",x"F1",x"C3",x"87",x"1F",x"01",x"FF",x"7C",x"C6",x"0E",x"3C",x"78",x"E0",x"FE",x"00",x"81",x"F3",x"E7",x"C3",x"F9",x"39",x"83",x"FF",x"7E",x"0C",x"18",x"3C",x"06",x"C6",x"7C",x"00",
																	x"E3",x"C3",x"93",x"33",x"01",x"F3",x"F3",x"FF",x"1C",x"3C",x"6C",x"CC",x"FE",x"0C",x"0C",x"00",x"03",x"3F",x"03",x"F9",x"F9",x"39",x"83",x"FF",x"FC",x"C0",x"FC",x"06",x"06",x"C6",x"7C",x"00",x"C3",x"9F",x"3F",x"03",x"39",x"39",x"83",x"FF",x"3C",x"60",x"C0",x"FC",x"C6",x"C6",x"7C",x"00",x"01",x"39",x"F3",x"E7",x"CF",x"CF",x"CF",x"FF",x"FE",x"C6",x"0C",x"18",x"30",x"30",x"30",x"00",
																	x"83",x"39",x"39",x"83",x"39",x"39",x"83",x"FF",x"7C",x"C6",x"C6",x"7C",x"C6",x"C6",x"7C",x"00",x"83",x"39",x"39",x"81",x"F9",x"F3",x"87",x"FF",x"7C",x"C6",x"C6",x"7E",x"06",x"0C",x"78",x"00",x"C7",x"93",x"39",x"39",x"01",x"39",x"39",x"FF",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"03",x"39",x"39",x"03",x"39",x"39",x"03",x"FF",x"FC",x"C6",x"C6",x"FC",x"C6",x"C6",x"FC",x"00",
																	x"C3",x"99",x"3F",x"3F",x"3F",x"99",x"C3",x"FF",x"3C",x"66",x"C0",x"C0",x"C0",x"66",x"3C",x"00",x"07",x"33",x"39",x"39",x"39",x"33",x"07",x"FF",x"F8",x"CC",x"C6",x"C6",x"C6",x"CC",x"F8",x"00",x"01",x"3F",x"3F",x"03",x"3F",x"3F",x"01",x"FF",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"FE",x"00",x"01",x"3F",x"3F",x"03",x"3F",x"3F",x"3F",x"FF",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"C0",x"00",
																	x"C1",x"9F",x"3F",x"31",x"39",x"99",x"C1",x"FF",x"3E",x"60",x"C0",x"CE",x"C6",x"66",x"3E",x"00",x"39",x"39",x"39",x"01",x"39",x"39",x"39",x"FF",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"00",x"81",x"E7",x"E7",x"E7",x"E7",x"E7",x"81",x"FF",x"7E",x"18",x"18",x"18",x"18",x"18",x"7E",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
																	x"39",x"33",x"27",x"0F",x"07",x"23",x"31",x"FF",x"C6",x"CC",x"D8",x"F0",x"F8",x"DC",x"CE",x"00",x"9F",x"9F",x"9F",x"9F",x"9F",x"9F",x"81",x"FF",x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00",x"39",x"11",x"01",x"01",x"29",x"39",x"39",x"FF",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"00",x"39",x"19",x"09",x"01",x"21",x"31",x"39",x"FF",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"00",
																	x"83",x"39",x"39",x"39",x"39",x"39",x"83",x"FF",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"03",x"39",x"39",x"39",x"03",x"3F",x"3F",x"FF",x"FC",x"C6",x"C6",x"C6",x"FC",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"00",x"00",x"00",x"C0",x"60",x"30",x"10",x"10",x"03",x"39",x"39",x"31",x"07",x"23",x"31",x"FF",x"FC",x"C6",x"C6",x"CE",x"F8",x"DC",x"CE",x"00",
																	x"87",x"33",x"3F",x"83",x"F9",x"39",x"83",x"FF",x"78",x"CC",x"C0",x"7C",x"06",x"C6",x"7C",x"00",x"81",x"E7",x"E7",x"E7",x"E7",x"E7",x"E7",x"FF",x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"39",x"39",x"39",x"39",x"39",x"39",x"83",x"FF",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"39",x"39",x"39",x"11",x"83",x"C7",x"EF",x"FF",x"C6",x"C6",x"C6",x"EE",x"7C",x"38",x"10",x"00",
																	x"39",x"39",x"29",x"01",x"01",x"11",x"39",x"FF",x"C6",x"C6",x"D6",x"FE",x"FE",x"EE",x"C6",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"99",x"99",x"81",x"C3",x"E7",x"E7",x"E7",x"FF",x"66",x"66",x"7E",x"3C",x"18",x"18",x"18",x"00",x"0F",x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"10",x"18",x"0C",x"07",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C3",x"BD",x"66",x"5E",x"5E",x"66",x"BD",x"C3",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C",x"FF",x"DF",x"CF",x"07",x"03",x"01",x"00",x"FF",x"00",x"20",x"30",x"F8",x"FC",x"FE",x"FF",x"00",x"FF",x"83",x"83",x"FF",x"83",x"83",x"FF",x"FF",x"00",x"7C",x"7C",x"00",x"7C",x"7C",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"04",x"18",x"30",x"1C",x"00",x"00",x"00",x"00",x"06",x"1F",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"EC",x"FE",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"38",x"70",x"70",x"38",x"FC",x"F8",x"7C",x"E6",x"3F",x"7F",x"7F",x"3F",x"FF",x"FF",x"7F",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"F8",x"F0",x"F8",x"F0",x"F8",x"01",x"07",x"0F",x"0C",x"1E",x"1F",x"0F",x"1F",x"01",x"07",x"0F",x"0F",x"1F",x"1F",x"0F",x"1F",x"C1",x"C0",x"E0",x"F0",x"60",x"C4",x"06",x"82",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"10",x"60",x"00",x"FC",x"FE",x"FC",x"FE",x"FE",x"FC",x"FE",x"FE",
																	x"3F",x"1F",x"0F",x"1F",x"3F",x"1F",x"3F",x"7F",x"3F",x"1F",x"0F",x"1F",x"3F",x"1F",x"3F",x"7F",x"C8",x"F8",x"F0",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"02",x"01",x"00",x"91",x"F3",x"FB",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"BF",x"42",x"C4",x"82",x"17",x"3E",x"FF",x"FF",x"BF",x"FE",x"FC",x"FE",x"FF",x"FE",x"FF",x"BF",x"DF",
																	x"7F",x"FF",x"FF",x"FF",x"EE",x"6E",x"76",x"30",x"7F",x"FF",x"7F",x"6F",x"77",x"B7",x"BB",x"DF",x"F6",x"F6",x"E4",x"E4",x"C4",x"40",x"40",x"00",x"BF",x"7F",x"7F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"9B",x"99",x"89",x"00",x"00",x"7D",x"7D",x"7D",x"FD",x"FE",x"FE",x"FF",x"FF",x"DE",x"DD",x"4C",x"A4",x"A4",x"80",x"80",x"00",x"EC",x"EE",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"10",x"14",x"14",x"08",x"08",x"08",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"08",x"0C",x"24",x"00",x"00",x"00",x"00",x"00",x"08",x"0C",x"24",x"00",x"00",x"00",x"00",x"00",x"01",x"22",x"62",x"00",x"00",x"00",x"00",x"00",x"02",x"24",x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"0C",
																	x"00",x"00",x"00",x"00",x"00",x"80",x"84",x"CC",x"00",x"00",x"00",x"00",x"00",x"80",x"84",x"CC",x"00",x"00",x"00",x"00",x"40",x"20",x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"30",x"00",x"00",x"00",x"00",x"00",x"40",x"51",x"51",x"00",x"00",x"00",x"00",x"01",x"01",x"02",x"82",x"00",x"00",x"00",x"80",x"80",x"80",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"33",x"31",x"31",x"10",x"10",x"00",x"00",x"00",x"DD",x"DE",x"DE",x"EF",x"EF",x"FF",x"FF",x"FF",x"80",x"80",x"80",x"80",x"04",x"04",x"04",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"40",x"80",x"80",x"88",x"88",x"08",x"08",x"08",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"22",x"22",x"12",x"12",x"12",x"10",x"10",x"10",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"08",x"08",x"08",x"08",x"04",x"04",x"04",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"10",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"E0",x"0F",x"00",x"00",x"00",x"00",x"00",x"1C",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E3",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"26",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D9",x"00",x"FF",
																	x"00",x"00",x"00",x"00",x"40",x"40",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"BF",x"1F",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"4C",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B3",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"C7",x"18",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FF",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FD",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"FB",x"E6",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FD",x"F9",x"F3",x"F3",x"00",x"40",x"48",x"08",x"22",x"26",x"4D",x"6F",x"C0",x"C0",x"E0",x"E0",x"E0",x"E0",x"A2",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"42",x"D4",
																	x"E2",x"62",x"22",x"20",x"20",x"00",x"00",x"00",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"2C",x"64",x"64",x"60",x"40",x"40",x"00",x"00",x"DE",x"9F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"9B",x"99",x"18",x"10",x"00",x"00",x"00",x"DD",x"ED",x"EF",x"EF",x"EF",x"FF",x"FF",x"FF",x"17",x"06",x"06",x"06",x"04",x"04",x"00",x"00",x"FB",x"FB",x"FB",x"FB",x"FF",x"FF",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"01",x"1D",x"3F",x"1F",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"19",x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"01",x"80",x"80",x"60",x"F8",x"F8",x"F6",x"FF",x"FF",
																	x"03",x"02",x"06",x"07",x"01",x"02",x"07",x"06",x"03",x"03",x"07",x"07",x"01",x"03",x"07",x"06",x"00",x"00",x"00",x"80",x"00",x"00",x"C0",x"88",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"03",x"00",x"00",x"00",x"01",x"00",x"04",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"C0",x"60",x"E0",x"C0",x"80",x"C0",x"00",x"80",x"C0",x"E0",x"E0",x"C0",x"80",x"C0",
																	x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"90",x"F0",x"B9",x"7F",x"6F",x"0E",x"04",x"00",x"FF",x"FF",x"BF",x"7F",x"6F",x"0E",x"04",x"00",x"00",x"81",x"91",x"BB",x"EF",x"EF",x"66",x"26",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"46",x"00",x"03",x"02",x"8A",x"CF",x"7B",x"30",x"10",x"00",x"FF",x"FE",x"FE",x"FF",x"7B",x"30",x"10",x"00",
																	x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"16",x"1E",x"0E",x"0E",x"0F",x"0F",x"C7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"01",x"00",x"40",x"E0",x"E8",x"FC",x"FE",x"FF",x"FF",x"7F",x"3F",x"07",x"07",x"03",x"03",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"03",x"80",x"81",x"82",x"C3",x"C1",x"C0",x"C0",x"03",x"00",x"01",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"22",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"02",x"01",x"03",x"0E",x"04",x"06",x"1E",x"24",x"FE",x"FF",x"FF",x"FE",x"FC",x"FE",x"FE",x"F4",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"E0",x"E0",x"E0",x"E0",x"C0",x"20",x"00",x"80",x"00",x"00",x"06",x"1F",x"3F",x"DF",x"FF",x"7F",x"0F",x"07",x"06",x"06",x"03",x"04",x"00",x"00",x"0F",x"05",x"C0",x"D8",x"FC",x"FB",x"FF",x"FF",x"77",x"FF",x"FE",x"EC",x"80",x"00",x"00",x"00",x"FF",x"FF",x"DE",x"0C",x"00",x"00",x"80",x"80",x"70",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"F0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"02",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"03",x"1B",x"3F",x"DF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"BB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"02",x"01",x"40",x"21",x"61",x"10",x"18",x"01",x"83",x"01",x"C0",x"E1",x"E1",x"D0",x"F8",
																	x"00",x"00",x"80",x"00",x"20",x"E4",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"37",x"00",x"00",x"00",x"00",x"82",x"89",x"DE",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"76",x"00",x"00",x"00",x"40",x"80",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"80",x"00",x"00",x"00",x"03",x"00",x"01",x"02",x"03",x"01",x"00",x"00",x"03",x"00",x"01",x"03",x"03",x"01",x"00",x"00",
																	x"80",x"80",x"00",x"20",x"C0",x"88",x"79",x"6F",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"7F",x"6F",x"00",x"00",x"00",x"00",x"00",x"02",x"11",x"39",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"38",x"10",x"18",x"58",x"38",x"20",x"F0",x"A0",x"F8",x"F0",x"F8",x"F8",x"F8",x"E0",x"F0",x"A0",x"7B",x"79",x"79",x"7B",x"7B",x"7B",x"7F",x"7F",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"E0",x"C0",x"C0",x"C0",x"C0",x"80",x"80",x"80",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"EF",x"E5",x"39",x"0F",x"03",x"00",x"00",x"FE",x"EE",x"C4",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"80",x"80",x"C0",x"C0",x"E0",x"E0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"7F",x"7F",x"7F",x"7F",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"70",x"78",x"38",x"3C",x"1E",x"1F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"7E",x"7E",x"FE",x"FE",x"FF",x"FF",x"FF",x"00",x"20",x"20",x"00",x"40",x"40",x"00",x"00",x"90",x"F0",x"B9",x"7F",x"6F",x"0F",x"1F",x"3E",x"FF",x"FF",x"BF",x"7F",x"6F",x"0E",x"04",x"00",
																	x"00",x"81",x"91",x"BB",x"EF",x"EF",x"46",x"00",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"46",x"00",x"07",x"07",x"03",x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"40",x"40",x"00",x"10",x"00",x"00",x"01",x"03",x"07",x"0F",x"9F",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"78",x"F0",x"FC",x"FF",x"E0",x"C0",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"10",x"00",x"20",x"20",x"00",x"00",x"00",x"08",x"FF",x"FE",x"FE",x"FC",x"F8",x"F8",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"00",x"20",x"20",x"00",x"00",x"00",x"10",x"10",
																	x"F0",x"E0",x"E0",x"C0",x"C0",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"FE",x"CE",x"CE",x"E7",x"77",x"73",x"73",x"66",x"EE",x"56",x"56",x"7B",x"FB",x"BD",x"BD",x"E5",x"C7",x"C7",x"C6",x"C6",x"C4",x"84",x"84",x"E9",x"DB",x"DB",x"FB",x"FF",x"FF",x"FF",x"FF",x"2E",x"46",x"4F",x"4F",x"4F",x"5E",x"4C",x"08",x"4E",x"86",x"87",x"D7",x"F7",x"EF",x"FF",x"FF",
																	x"DD",x"7D",x"6F",x"66",x"B6",x"B2",x"90",x"90",x"CD",x"6D",x"77",x"FB",x"FB",x"FF",x"FF",x"FF",x"08",x"00",x"20",x"62",x"22",x"20",x"00",x"00",x"90",x"99",x"BD",x"FF",x"FF",x"FF",x"FF",x"FF",x"11",x"10",x"08",x"08",x"01",x"01",x"41",x"41",x"A2",x"A7",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"20",x"A8",x"88",x"84",x"0A",x"02",x"00",x"00",x"01",x"C1",x"E1",x"E9",x"FF",x"FF",x"FF",x"FF",
																	x"08",x"84",x"84",x"60",x"20",x"20",x"10",x"10",x"31",x"19",x"19",x"BD",x"FF",x"FF",x"FF",x"FF",x"01",x"03",x"05",x"07",x"0B",x"1F",x"37",x"3B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"80",x"80",x"E0",x"D0",x"F0",x"F0",x"F8",x"EC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"03",x"06",x"0B",x"1F",x"1D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"C0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"2F",x"7F",x"3D",x"DF",x"F7",x"7F",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"F8",x"F4",x"FE",x"FE",x"FC",x"FE",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0B",x"1F",x"2F",x"3F",x"5B",x"EF",x"FE",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"E0",x"D0",x"F8",x"F0",x"F8",x"F4",x"FC",x"EE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"EF",x"FF",x"7F",x"5B",x"2F",x"3B",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"EE",x"FA",x"FC",x"F4",x"F8",x"EC",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"5F",x"F7",x"7F",x"3F",x"6F",x"5B",x"3E",x"17",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"FE",x"F4",x"F8",x"FC",x"B4",x"D8",x"F8",x"D0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"E0",x"80",x"80",x"80",x"80",x"80",x"80",x"C0",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"E0",x"C0",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"FF",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
																	x"08",x"0C",x"14",x"3E",x"5E",x"7D",x"3E",x"5F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"10",x"38",x"5C",x"7C",x"FA",x"5E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3D",x"2E",x"7E",x"2C",x"08",x"08",x"08",x"08",x"FF",x"FF",x"FF",x"FF",x"F7",x"F7",x"F7",x"F7",x"FF",x"ED",x"BE",x"7C",x"38",x"10",x"10",x"10",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"EF",x"EF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"0F",x"0F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"0F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"60",x"38",x"0E",x"0F",x"1F",x"03",x"01",x"00",x"E0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"0F",x"3F",x"7F",x"7F",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"1F",x"3F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"EF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"3F",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"1F",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"18",x"0C",x"07",x"07",x"0F",x"1F",x"03",x"00",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"80",x"F0",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"80",x"F0",x"FC",x"FE",x"FF",x"80",x"F0",x"F8",x"FE",x"FF",x"0F",x"03",x"00",x"80",x"F0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"F0",x"FC",x"FF",x"FF",x"00",x"00",x"00",x"00",x"F0",x"FC",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"FF",x"7F",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"E0",x"38",x"0F",x"07",x"07",x"0F",x"03",x"00",x"E0",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"E0",x"F0",x"F8",x"FF",x"FF",x"00",x"00",x"00",x"E0",x"F0",x"F8",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"FE",x"1F",x"07",x"07",x"0F",x"1F",x"03",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FF",x"00",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FF",x"03",x"01",x"03",x"1F",x"0F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"07",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"80",x"F0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"80",x"F0",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"FE",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"1F",x"FF",x"3F",x"1F",x"07",x"07",x"0F",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"80",x"E0",x"F0",x"FC",x"FF",x"FF",x"FF",x"FF",x"80",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"3F",x"1F",x"1F",x"1F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"C0",x"F0",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"01",x"51",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"12",x"52",x"00",x"00",x"00",x"00",x"10",x"22",x"2B",x"9B",x"00",x"00",x"00",x"00",x"00",x"02",x"49",x"DD",x"FF",x"FF",x"DF",x"BF",x"BF",x"FF",x"FF",x"FF",x"00",x"38",x"7C",x"FE",x"FE",x"FE",x"7C",x"38",
																	x"FF",x"C7",x"83",x"01",x"01",x"01",x"83",x"C7",x"00",x"38",x"7C",x"FE",x"FE",x"FE",x"7C",x"38",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"70",x"F0",x"30",x"76",x"FE",x"FC",x"78",x"FF",x"8F",x"0F",x"CF",x"89",x"01",x"03",x"87",x"00",x"70",x"F0",x"30",x"76",x"FE",x"FC",x"78",x"FF",x"FF",x"55",x"55",x"55",x"55",x"55",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"FF",x"EF",x"EF",x"EF",x"EF",x"FF",x"EF",x"FF",x"18",x"2C",x"2C",x"2C",x"2C",x"00",x"2C",x"00",x"FF",x"84",x"9C",x"84",x"E4",x"E4",x"84",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"90",x"92",x"12",x"92",x"92",x"90",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"FF",x"43",x"67",x"67",x"67",x"67",x"67",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"FF",x"3F",x"9F",x"CF",x"E7",x"F3",x"F9",x"FC",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
																	x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"FF",x"FC",x"F9",x"F3",x"E7",x"CF",x"9F",x"3F",x"7F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"F9",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
																	x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BF",x"BF",x"BF",x"BF",x"BF",x"BF",x"BF",x"BF",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",
																	x"F9",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"1F",x"FF",x"FF",x"FF",x"FF",
																	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"1F",x"1F",x"0F",x"0F",x"1F",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"93",x"93",x"F7",x"FF",x"00",x"00",x"00",x"00",x"6C",x"6C",x"08",x"00",x"FF",x"FF",x"FF",x"FF",x"9F",x"9F",x"FF",x"FF",x"00",x"00",x"00",x"00",x"60",x"60",x"00",x"00",
																	x"E0",x"F8",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FE",x"FE",x"FC",x"F8",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"1F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"7F",x"7F",x"3F",x"1F",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"C3",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C3",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"00",x"00",x"01",x"01",x"03",x"03",x"07",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"07",x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
																	x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"10",x"30",x"60",x"C0",x"00",x"00",x"00",x"00",x"99",x"99",x"99",x"BB",x"FF",x"33",x"33",x"FF",x"66",x"66",x"66",x"44",x"00",x"CC",x"CC",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"0F",x"00",x"00",x"00",x"07",x"0C",x"18",x"10",x"10");
	
	
	constant DONKEY_KONG_CHR_ROM : CHR_ROM_ARRAY := (x"00",x"03",x"07",x"07",x"09",x"09",x"1C",x"00",x"00",x"03",x"07",x"00",x"06",x"06",x"03",x"03",x"0F",x"0F",x"0F",x"FF",x"FF",x"FC",x"81",x"01",x"00",x"10",x"3C",x"3F",x"3F",x"3C",x"00",x"00",x"00",x"C0",x"F8",x"80",x"20",x"90",x"3C",x"00",x"00",x"C0",x"F8",x"60",x"DC",x"6E",x"C0",x"F8",x"C0",x"C0",x"C0",x"F0",x"F0",x"E0",x"C0",x"E0",x"50",x"38",x"30",x"F0",x"F0",x"E0",x"00",x"00",x"07",x"0F",x"0F",x"12",x"13",x"38",x"00",x"0F",x"07",x"0F",x"00",x"0D",x"0C",x"07",x"07",x"00",x"1F",x"1F",x"1F",x"18",x"19",x"1E",x"1C",x"1E",x"01",x"03",x"01",x"17",x"1F",x"1E",x"00",x"00",x"80",x"F0",x"00",x"40",x"20",x"78",x"00",x"C0",x"80",x"F0",x"C0",x"B8",x"DC",x"80",x"F0",x"00",x"E0",x"60",x"F0",x"F0",x"F0",x"E0",x"E0",x"F0",x"80",x"E0",x"F0",x"F0",x"F0",x"E0",x"00",x"00",
															x"07",x"0F",x"0F",x"12",x"13",x"38",x"00",x"3F",x"07",x"0F",x"00",x"0D",x"0C",x"07",x"07",x"03",x"3F",x"0E",x"0F",x"1F",x"3F",x"7C",x"70",x"38",x"C3",x"E3",x"CF",x"1F",x"3F",x"0C",x"00",x"00",x"80",x"F0",x"00",x"40",x"20",x"78",x"00",x"C0",x"80",x"F0",x"C0",x"B8",x"DC",x"80",x"F0",x"06",x"F0",x"F8",x"E4",x"FC",x"FC",x"7C",x"00",x"00",x"8E",x"E6",x"E0",x"F0",x"F0",x"70",x"00",x"00",x"00",x"02",x"06",x"07",x"09",x"09",x"1D",x"03",x"01",x"03",x"07",x"00",x"06",x"06",x"02",x"00",x"0F",x"0F",x"0F",x"FF",x"FF",x"FC",x"81",x"01",x"00",x"00",x"0C",x"3F",x"3F",x"3C",x"00",x"00",x"00",x"00",x"38",x"C0",x"E0",x"D0",x"FC",x"C0",x"C0",x"C0",x"F8",x"20",x"1C",x"2E",x"00",x"38",x"E0",x"E0",x"B0",x"F0",x"F0",x"E0",x"C0",x"E0",x"00",x"60",x"F0",x"F0",x"F0",x"E0",x"00",x"00",
															x"00",x"03",x"07",x"07",x"09",x"09",x"1C",x"00",x"00",x"03",x"07",x"00",x"06",x"06",x"03",x"03",x"0F",x"0F",x"0F",x"FF",x"FF",x"FC",x"81",x"01",x"00",x"00",x"0C",x"3F",x"3F",x"3C",x"00",x"00",x"00",x"C0",x"F8",x"80",x"20",x"90",x"3C",x"00",x"00",x"C0",x"F8",x"60",x"DC",x"6E",x"C0",x"F8",x"E0",x"F0",x"F0",x"F0",x"F0",x"E0",x"C0",x"E0",x"47",x"0F",x"0E",x"F0",x"F0",x"E0",x"00",x"00",x"04",x"0C",x"0C",x"13",x"13",x"3B",x"07",x"0F",x"07",x"0F",x"03",x"0C",x"0C",x"04",x"00",x"00",x"0F",x"0F",x"0F",x"1F",x"1F",x"1E",x"1C",x"1E",x"00",x"01",x"0F",x"1F",x"1F",x"1E",x"00",x"00",x"00",x"70",x"00",x"C0",x"A0",x"F8",x"80",x"C0",x"80",x"F0",x"C0",x"38",x"5C",x"00",x"70",x"40",x"E0",x"60",x"F0",x"F0",x"F0",x"E0",x"E0",x"F0",x"C0",x"E0",x"F0",x"F0",x"F0",x"E0",x"00",x"00",
															x"07",x"0F",x"0F",x"12",x"13",x"38",x"00",x"0F",x"07",x"0F",x"00",x"0D",x"0C",x"07",x"07",x"01",x"1F",x"1F",x"1F",x"1F",x"1F",x"1E",x"1C",x"1E",x"00",x"00",x"13",x"1F",x"1F",x"1E",x"00",x"00",x"80",x"F0",x"00",x"40",x"20",x"78",x"00",x"C0",x"80",x"F0",x"C0",x"B8",x"DC",x"80",x"F0",x"80",x"F8",x"F8",x"F0",x"F0",x"F0",x"E0",x"E0",x"F0",x"07",x"07",x"FE",x"F0",x"F0",x"E0",x"00",x"00",x"04",x"0C",x"0C",x"13",x"13",x"3F",x"07",x"0F",x"07",x"0F",x"03",x"0C",x"0C",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"1F",x"3F",x"7C",x"70",x"38",x"01",x"01",x"0F",x"1F",x"3F",x"1C",x"00",x"00",x"00",x"70",x"00",x"C0",x"A0",x"F8",x"80",x"C0",x"80",x"F0",x"C0",x"38",x"5C",x"00",x"70",x"40",x"C0",x"60",x"E4",x"FC",x"FC",x"7C",x"00",x"00",x"C0",x"E0",x"E0",x"F0",x"F0",x"70",x"00",x"00",
															x"07",x"0F",x"0F",x"12",x"13",x"38",x"00",x"07",x"07",x"0F",x"00",x"0D",x"0C",x"07",x"07",x"01",x"0F",x"0F",x"0F",x"1F",x"3F",x"7C",x"70",x"38",x"00",x"00",x"09",x"1F",x"3F",x"1C",x"00",x"00",x"80",x"F0",x"00",x"40",x"20",x"78",x"00",x"C0",x"80",x"F0",x"C0",x"B8",x"DC",x"80",x"F0",x"80",x"F8",x"F8",x"E0",x"FC",x"FC",x"7C",x"00",x"00",x"07",x"07",x"EE",x"F0",x"F0",x"70",x"00",x"00",x"00",x"07",x"07",x"0F",x"0F",x"38",x"7F",x"7F",x"00",x"07",x"03",x"00",x"00",x"07",x"04",x"04",x"1F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"07",x"1E",x"1F",x"1F",x"1F",x"0F",x"08",x"00",x"00",x"00",x"E0",x"F8",x"FC",x"FC",x"1C",x"F8",x"F8",x"38",x"F8",x"C0",x"00",x"00",x"E0",x"20",x"20",x"F8",x"FC",x"FC",x"F8",x"78",x"80",x"C0",x"C0",x"78",x"FC",x"FC",x"F8",x"00",x"80",x"00",x"00",
															x"00",x"03",x"07",x"07",x"09",x"09",x"1C",x"00",x"00",x"03",x"07",x"00",x"06",x"06",x"03",x"63",x"1F",x"0F",x"07",x"37",x"7F",x"DF",x"0F",x"06",x"E0",x"21",x"01",x"07",x"07",x"1F",x"0F",x"06",x"00",x"C0",x"F8",x"80",x"20",x"90",x"3C",x"00",x"00",x"C0",x"F8",x"60",x"DC",x"6E",x"C0",x"FB",x"E4",x"FE",x"70",x"F1",x"FF",x"FF",x"00",x"00",x"83",x"C0",x"F0",x"F0",x"FC",x"FC",x"00",x"00",x"07",x"0F",x"0F",x"12",x"13",x"38",x"70",x"FF",x"07",x"0F",x"00",x"0D",x"0C",x"07",x"0F",x"02",x"DF",x"1E",x"1F",x"1F",x"1F",x"0F",x"07",x"01",x"01",x"F3",x"5F",x"1F",x"1F",x"4F",x"37",x"C0",x"80",x"F0",x"00",x"40",x"20",x"78",x"00",x"FC",x"80",x"F0",x"C0",x"B8",x"DC",x"80",x"F0",x"00",x"F0",x"E0",x"E0",x"F0",x"FA",x"FE",x"FC",x"D8",x"8F",x"E7",x"E0",x"F0",x"C8",x"88",x"10",x"00",
															x"00",x"00",x"07",x"08",x"10",x"20",x"40",x"40",x"00",x"00",x"00",x"07",x"08",x"10",x"20",x"20",x"40",x"40",x"20",x"10",x"08",x"07",x"00",x"00",x"20",x"20",x"10",x"08",x"07",x"00",x"00",x"00",x"00",x"00",x"E0",x"10",x"08",x"04",x"02",x"02",x"00",x"00",x"00",x"E0",x"10",x"08",x"04",x"04",x"02",x"02",x"04",x"08",x"10",x"E0",x"00",x"00",x"04",x"04",x"08",x"10",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"04",x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"03",x"04",x"08",x"10",x"08",x"04",x"03",x"00",x"00",x"00",x"00",x"08",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"20",x"10",x"08",x"00",x"00",x"00",x"00",x"00",x"C0",x"20",x"10",x"08",x"10",x"20",x"C0",x"00",x"00",x"00",x"00",x"10",x"20",x"C0",x"00",x"00",x"00",x"00",x"00",
															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"21",x"10",x"00",x"00",x"00",x"01",x"01",x"40",x"00",x"00",x"00",x"00",x"60",x"00",x"00",x"10",x"21",x"01",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"40",x"01",x"01",x"00",x"00",x"00",x"00",x"08",x"10",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"0C",x"00",x"00",x"10",x"08",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"04",x"00",x"00",
															x"04",x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"0F",x"07",x"03",x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"42",x"39",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"0F",x"1F",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"1F",x"FF",x"FF",x"FF",x"F8",x"F7",x"EF",x"FF",x"FF",x"FE",x"7E",x"3E",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",
															x"00",x"00",x"00",x"C0",x"E0",x"F0",x"DB",x"F6",x"00",x"80",x"80",x"C0",x"E0",x"F0",x"FF",x"FF",x"CB",x"E0",x"C4",x"02",x"D1",x"E1",x"D1",x"83",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"FF",x"E0",x"8F",x"6E",x"44",x"EE",x"60",x"FF",x"FF",x"FF",x"F0",x"80",x"00",x"00",x"9F",x"83",x"E0",x"E4",x"C6",x"61",x"33",x"1F",x"0F",x"FF",x"FF",x"F9",x"F9",x"7F",x"3F",x"1F",x"0F",x"00",x"00",x"00",x"03",x"07",x"0F",x"5B",x"A7",x"00",x"01",x"01",x"03",x"07",x"0F",x"FF",x"FF",x"73",x"07",x"27",x"40",x"8B",x"87",x"8B",x"C1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"FF",x"0F",x"E1",x"EC",x"44",x"EE",x"0C",x"FF",x"FF",x"FF",x"1F",x"03",x"01",x"01",x"F3",x"80",x"0E",x"4E",x"C6",x"0C",x"98",x"F0",x"E0",x"FF",x"FF",x"3F",x"3F",x"FC",x"F8",x"F0",x"E0",
															x"00",x"42",x"9C",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"F8",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",x"F8",x"FF",x"FF",x"FF",x"1F",x"EF",x"F7",x"FF",x"FF",x"FE",x"7C",x"70",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"80",x"00",x"00",x"00",x"00",x"00",x"F0",x"E0",x"C0",x"00",x"00",x"80",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"00",x"00",x"1F",x"3F",x"3F",x"7F",x"7F",x"7F",x"00",x"0F",x"28",x"5C",x"3F",x"7F",x"7F",x"7F",x"7F",x"3E",x"1F",x"1F",x"0F",x"0F",x"0F",x"07",x"7F",x"3E",x"1F",x"1F",x"08",x"00",x"00",x"00",x"00",x"60",x"F0",x"F8",x"F8",x"F8",x"FC",x"FC",x"00",x"80",x"40",x"C4",x"F6",x"FE",x"FC",x"FC",x"F8",x"F0",x"F0",x"E0",x"80",x"80",x"C0",x"C0",x"F8",x"F0",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"1F",x"3F",x"7F",x"FF",x"FF",x"3E",x"0F",x"00",x"1C",x"3F",x"7F",x"FF",x"FF",x"3E",x"70",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"F0",x"FC",x"FE",x"FE",x"FF",x"FC",x"00",x"60",x"F0",x"F8",x"FC",x"FC",x"FC",x"FF",x"7C",x"FC",x"F8",x"F0",x"E0",x"00",x"00",x"00",x"7C",x"FC",x"88",x"00",x"00",x"00",x"00",x"00",
															x"00",x"07",x"07",x"0F",x"0F",x"00",x"1F",x"3F",x"00",x"07",x"03",x"00",x"00",x"07",x"04",x"04",x"7F",x"7F",x"1F",x"1F",x"1F",x"1E",x"0F",x"1F",x"0C",x"9E",x"FF",x"1F",x"1F",x"1E",x"0F",x"00",x"00",x"E0",x"E0",x"F0",x"F0",x"00",x"F8",x"FC",x"00",x"E0",x"C0",x"00",x"00",x"E0",x"20",x"20",x"FE",x"FE",x"F8",x"F8",x"F8",x"78",x"F0",x"F8",x"30",x"79",x"FF",x"F8",x"F8",x"78",x"F0",x"00",x"03",x"07",x"05",x"08",x"1B",x"19",x"05",x"3F",x"03",x"07",x"02",x"07",x"04",x"46",x"E3",x"C2",x"3F",x"0F",x"05",x"37",x"3F",x"3F",x"3E",x"1C",x"42",x"07",x"07",x"07",x"07",x"03",x"02",x"00",x"E0",x"F0",x"50",x"08",x"6C",x"CC",x"D0",x"FE",x"E0",x"F0",x"A0",x"F0",x"90",x"32",x"E3",x"21",x"FE",x"F8",x"D0",x"FB",x"FF",x"FF",x"3E",x"0C",x"20",x"70",x"F0",x"F8",x"F8",x"F0",x"30",x"00",
															x"00",x"00",x"79",x"F9",x"F3",x"FF",x"7B",x"3F",x"00",x"01",x"00",x"00",x"00",x"1E",x"7F",x"3E",x"3F",x"3F",x"7B",x"7F",x"FB",x"F1",x"79",x"38",x"3C",x"3E",x"7F",x"7E",x"18",x"00",x"00",x"00",x"00",x"00",x"80",x"B0",x"B8",x"C6",x"93",x"F7",x"C0",x"E0",x"40",x"00",x"00",x"3A",x"EF",x"4B",x"E3",x"F7",x"93",x"C6",x"B8",x"B0",x"80",x"00",x"5F",x"4B",x"EF",x"3A",x"00",x"00",x"60",x"C0",x"30",x"7C",x"FF",x"FF",x"DF",x"0B",x"1F",x"7F",x"00",x"0C",x"0F",x"1F",x"1F",x"0F",x"0E",x"04",x"7F",x"0B",x"33",x"36",x"10",x"0A",x"0F",x"07",x"84",x"C7",x"4C",x"09",x"0F",x"05",x"0F",x"07",x"38",x"7C",x"FC",x"FC",x"EC",x"A0",x"F0",x"FC",x"00",x"40",x"C0",x"E0",x"E0",x"E0",x"E0",x"42",x"FC",x"A0",x"98",x"D8",x"10",x"A0",x"E0",x"C0",x"43",x"C7",x"62",x"20",x"E0",x"40",x"E0",x"C0",
															x"00",x"01",x"0D",x"1D",x"63",x"C9",x"EF",x"C7",x"03",x"04",x"00",x"00",x"5C",x"F7",x"D2",x"FA",x"EF",x"C9",x"63",x"1D",x"0D",x"01",x"00",x"00",x"D2",x"F7",x"5C",x"00",x"00",x"02",x"07",x"03",x"1C",x"9E",x"8F",x"DF",x"FE",x"DE",x"FC",x"FC",x"00",x"00",x"00",x"18",x"7E",x"FE",x"7C",x"3C",x"FC",x"DE",x"FF",x"CF",x"9F",x"9E",x"00",x"00",x"7C",x"FE",x"78",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"00",x"00",x"1E",x"3F",x"7D",x"78",x"00",x"00",x"01",x"00",x"00",x"20",x"7C",x"78",x"7C",x"FB",x"FF",x"FF",x"5F",x"1F",x"1F",x"1F",x"7C",x"FE",x"FF",x"FE",x"7C",x"60",x"E0",x"E1",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"00",x"7C",x"82",x"01",x"82",x"7C",x"00",x"00",x"00",x"00",x"21",x"A2",x"A3",x"B3",x"8F",x"27",x"FE",x"10",x"19",x"5A",x"DF",x"4F",x"73",x"DB",x"02",
															x"00",x"00",x"00",x"00",x"03",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"03",x"0C",x"10",x"22",x"20",x"1F",x"1F",x"0F",x"03",x"00",x"00",x"00",x"00",x"21",x"23",x"10",x"0C",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"F8",x"00",x"00",x"00",x"C0",x"30",x"08",x"64",x"C4",x"F8",x"F8",x"F0",x"C0",x"00",x"00",x"00",x"00",x"84",x"04",x"08",x"30",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"03",x"0C",x"10",x"26",x"23",x"1F",x"1F",x"0F",x"03",x"00",x"00",x"00",x"00",x"21",x"20",x"10",x"0C",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"F8",x"00",x"00",x"00",x"C0",x"30",x"08",x"44",x"04",x"F8",x"F8",x"F0",x"C0",x"00",x"00",x"00",x"00",x"84",x"C4",x"08",x"30",x"C0",x"00",x"00",x"00",
															x"00",x"00",x"00",x"00",x"03",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"03",x"0C",x"10",x"20",x"21",x"1F",x"1F",x"0F",x"03",x"00",x"00",x"00",x"00",x"23",x"26",x"10",x"0C",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"F8",x"00",x"00",x"00",x"C0",x"30",x"08",x"C4",x"84",x"F8",x"F8",x"F0",x"C0",x"00",x"00",x"00",x"00",x"04",x"44",x"08",x"30",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"03",x"0C",x"10",x"23",x"21",x"1F",x"1F",x"0F",x"03",x"00",x"00",x"00",x"00",x"20",x"22",x"10",x"0C",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"F8",x"F8",x"00",x"00",x"00",x"C0",x"30",x"08",x"04",x"84",x"F8",x"F8",x"F0",x"C0",x"00",x"00",x"00",x"00",x"C4",x"64",x"08",x"30",x"C0",x"00",x"00",x"00",
															x"00",x"00",x"00",x"0F",x"30",x"60",x"3F",x"7F",x"00",x"00",x"00",x"00",x"2F",x"3F",x"60",x"20",x"7F",x"3F",x"60",x"30",x"0F",x"00",x"00",x"00",x"20",x"60",x"3F",x"2F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"06",x"03",x"FE",x"FF",x"00",x"00",x"00",x"00",x"FA",x"FE",x"03",x"02",x"FF",x"FE",x"03",x"06",x"F8",x"00",x"00",x"00",x"02",x"03",x"FE",x"FA",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2F",x"3F",x"60",x"20",x"00",x"00",x"00",x"0F",x"30",x"60",x"3F",x"7F",x"20",x"60",x"3F",x"2F",x"00",x"00",x"00",x"00",x"7F",x"3F",x"60",x"30",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FA",x"FE",x"03",x"02",x"00",x"00",x"00",x"F8",x"06",x"03",x"FE",x"FF",x"02",x"03",x"FE",x"FA",x"00",x"00",x"00",x"00",x"FF",x"FE",x"03",x"06",x"F8",x"00",x"00",x"00",
															x"00",x"44",x"00",x"41",x"20",x"4B",x"27",x"1F",x"00",x"00",x"00",x"40",x"20",x"00",x"00",x"01",x"0F",x"1E",x"1F",x"1F",x"1F",x"0F",x"0F",x"03",x"03",x"07",x"06",x"06",x"07",x"03",x"00",x"00",x"00",x"20",x"50",x"20",x"60",x"48",x"E0",x"F0",x"00",x"00",x"40",x"00",x"00",x"08",x"00",x"40",x"F8",x"78",x"3C",x"3C",x"3C",x"FC",x"F8",x"E0",x"E0",x"F0",x"D0",x"D0",x"F0",x"E0",x"00",x"00",x"10",x"01",x"2A",x"0C",x"A6",x"17",x"1F",x"1F",x"00",x"00",x"02",x"00",x"80",x"00",x"03",x"07",x"5E",x"3C",x"3D",x"3D",x"3E",x"1F",x"0F",x"07",x"07",x"0F",x"0E",x"0E",x"0F",x"07",x"03",x"00",x"00",x"00",x"80",x"C8",x"60",x"E0",x"F4",x"F8",x"00",x"00",x"00",x"08",x"00",x"80",x"24",x"C0",x"7C",x"1C",x"2E",x"2E",x"1E",x"FC",x"F8",x"E0",x"F0",x"F8",x"D8",x"D8",x"F8",x"F0",x"C0",x"00",
															x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"92",x"54",x"38",x"FE",x"38",x"54",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"00",x"00",x"00",x"00",x"00",x"23",x"97",x"2F",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"6E",x"EF",x"F7",x"FF",x"7F",x"3F",x"5F",x"0F",x"07",x"07",x"03",x"27",x"1F",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"FE",x"5E",x"00",x"00",x"00",x"00",x"00",x"F0",x"F8",x"AC",x"5E",x"0C",x"9E",x"FE",x"FE",x"FE",x"F8",x"C0",x"AC",x"F8",x"F8",x"F8",x"F0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"2F",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"4E",x"6E",x"FE",x"7F",x"3F",x"1F",x"0F",x"03",x"07",x"07",x"07",x"27",x"1F",x"07",x"01",x"00",x"00",x"00",x"00",x"00",x"F8",x"FC",x"FE",x"56",x"00",x"00",x"00",x"00",x"00",x"F0",x"F8",x"AC",x"56",x"0C",x"0E",x"1F",x"FF",x"FF",x"FE",x"F8",x"AC",x"F8",x"F8",x"FC",x"FC",x"F8",x"F0",x"00",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"00",x"07",x"08",x"10",x"10",x"20",x"20",x"20",x"00",x"07",x"08",x"10",x"10",x"20",x"20",x"20",x"1F",x"2F",x"37",x"3A",x"3D",x"3E",x"3F",x"00",x"1F",x"3F",x"3F",x"3F",x"3E",x"3F",x"3F",x"00",x"00",x"05",x"19",x"33",x"63",x"C7",x"C7",x"C4",x"00",x"07",x"1F",x"3F",x"7F",x"FF",x"FF",x"DD",x"80",x"00",x"00",x"00",x"00",x"03",x"03",x"00",x"89",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"07",x"00",x"00",x"0F",x"00",x"80",x"63",x"1E",x"00",x"0F",x"0F",x"00",x"1F",x"7F",x"1C",x"00",x"00",x"01",x"03",x"19",x"3C",x"19",x"23",x"51",x"20",x"01",x"02",x"19",x"24",x"19",x"22",x"11",x"2C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"07",x"03",x"03",x"01",x"01",x"01",x"00",
															x"00",x"3F",x"1F",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0D",x"19",x"11",x"00",x"01",x"00",x"01",x"00",x"1F",x"3F",x"29",x"19",x"0D",x"07",x"03",x"01",x"00",x"00",x"00",x"FC",x"F8",x"00",x"80",x"00",x"80",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"B0",x"98",x"88",x"00",x"80",x"00",x"80",x"00",x"F8",x"FC",x"94",x"98",x"B0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"41",x"01",x"01",x"00",x"1F",x"3F",x"0F",x"79",x"A1",x"79",x"0F",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"82",x"80",x"80",x"00",x"F8",x"FC",x"F0",x"9E",x"85",x"9E",x"F0",x"80",x"00",x"00",
															x"00",x"00",x"00",x"1E",x"3F",x"3F",x"3F",x"3F",x"00",x"00",x"00",x"1E",x"3F",x"3F",x"3F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"1F",x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"7E",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"3C",x"7E",x"FE",x"FE",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"08",x"19",x"09",x"09",x"09",x"09",x"1C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"05",x"05",x"19",x"05",x"05",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"21",x"21",x"3D",x"05",x"05",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"25",x"25",x"19",x"25",x"25",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"29",x"29",x"29",x"29",x"29",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"63",x"31",x"1F",x"00",x"00",x"00",x"00",x"3C",x"B6",x"7C",x"F8",x"00",x"00",x"FC",x"FE",x"C0",x"40",x"80",x"00",x"03",x"03",x"03",x"07",x"0C",x"1B",x"77",x"07",x"7F",x"3F",x"53",x"07",x"0C",x"1B",x"07",x"07",
															x"0F",x"0F",x"1F",x"3F",x"7F",x"3F",x"00",x"00",x"0F",x"0F",x"03",x"38",x"3F",x"0E",x"1C",x"0E",x"E0",x"F0",x"F0",x"F0",x"18",x"FC",x"FC",x"FC",x"00",x"90",x"F0",x"F0",x"18",x"FC",x"F0",x"F8",x"F8",x"FC",x"FF",x"FF",x"FE",x"F0",x"00",x"00",x"F8",x"F0",x"87",x"3D",x"FE",x"1C",x"08",x"00",x"03",x"03",x"03",x"03",x"01",x"00",x"07",x"1F",x"7F",x"3F",x"53",x"03",x"01",x"00",x"07",x"1F",x"FF",x"FF",x"7F",x"3F",x"0F",x"03",x"00",x"00",x"CF",x"63",x"38",x"3E",x"7B",x"30",x"18",x"00",x"E0",x"F0",x"F0",x"E0",x"FE",x"3C",x"F0",x"FC",x"00",x"90",x"F0",x"E0",x"F8",x"38",x"F0",x"F0",x"FC",x"F8",x"F8",x"F8",x"F8",x"F8",x"F8",x"00",x"F8",x"F8",x"F8",x"38",x"80",x"F8",x"00",x"5C",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"03",x"33",x"19",x"0F",x"3F",x"1F",x"00",x"01",x"03",x"33",x"19",x"0F",x"3F",x"1F",x"2B",x"07",x"05",x"0D",x"0B",x"1B",x"1B",x"3B",x"2B",x"07",x"05",x"0D",x"0B",x"1B",x"1B",x"03",x"09",x"00",x"07",x"07",x"0F",x"0D",x"01",x"00",x"01",x"00",x"03",x"05",x"0E",x"0D",x"01",x"00",x"F8",x"FC",x"F8",x"EC",x"F8",x"F0",x"C0",x"C0",x"F8",x"FC",x"C0",x"40",x"80",x"80",x"00",x"80",
															x"F0",x"F8",x"F8",x"E8",x"CC",x"E6",x"FB",x"FF",x"D0",x"F8",x"F8",x"E8",x"CC",x"E6",x"F8",x"FE",x"FF",x"FE",x"FE",x"FE",x"FE",x"8F",x"00",x"00",x"FE",x"FE",x"06",x"F8",x"0E",x"80",x"00",x"00",x"01",x"0F",x"00",x"00",x"04",x"1E",x"00",x"03",x"01",x"0F",x"07",x"1D",x"3B",x"01",x"0F",x"02",x"07",x"0F",x"1F",x"0F",x"07",x"0F",x"0F",x"03",x"02",x"03",x"02",x"77",x"17",x"01",x"00",x"00",x"E0",x"F0",x"F0",x"48",x"C8",x"9C",x"00",x"F0",x"E0",x"F0",x"00",x"B0",x"30",x"60",x"F0",x"10",x"F8",x"FC",x"FC",x"F8",x"F8",x"78",x"70",x"60",x"30",x"F0",x"D0",x"FC",x"FE",x"08",x"00",x"00",x"00",x"00",x"7C",x"8A",x"FE",x"FE",x"FE",x"FE",x"00",x"10",x"00",x"74",x"00",x"00",x"00",x"00",x"FE",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",
															x"07",x"0B",x"0F",x"0B",x"0B",x"0B",x"0B",x"07",x"00",x"04",x"00",x"14",x"04",x"04",x"04",x"00",x"C0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"00",x"00",x"00",x"1F",x"00",x"00",x"00",x"00",x"03",x"07",x"07",x"07",x"07",x"07",x"07",x"03",x"00",x"00",x"00",x"F8",x"00",x"00",x"00",x"00",x"E0",x"D0",x"D0",x"D0",x"D0",x"F0",x"D0",x"E0",x"00",x"20",x"20",x"28",x"20",x"00",x"20",x"00",x"00",x"01",x"13",x"37",x"3B",x"74",x"7A",x"3E",x"00",x"00",x"08",x"25",x"12",x"53",x"33",x"39",x"D8",x"98",x"A8",x"D8",x"DA",x"74",x"28",x"C8",x"08",x"80",x"30",x"9C",x"CA",x"B8",x"98",x"78",x"08",x"59",x"30",x"71",x"79",x"2B",x"36",x"16",x"00",x"08",x"00",x"40",x"00",x"31",x"3D",x"19",x"C6",x"C4",x"CC",x"CC",x"B8",x"7C",x"EC",x"C8",x"00",x"80",x"C0",x"C0",x"C0",x"88",x"B8",x"B8",
															x"38",x"4C",x"C6",x"C6",x"C6",x"64",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"38",x"18",x"18",x"18",x"18",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"0E",x"3C",x"78",x"E0",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"0C",x"18",x"3C",x"06",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"3C",x"6C",x"CC",x"FE",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"C0",x"FC",x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"60",x"C0",x"FC",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"C6",x"0C",x"18",x"30",x"30",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"78",x"C4",x"E4",x"78",x"86",x"86",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"7E",x"06",x"0C",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"C6",x"C6",x"FC",x"C6",x"C6",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"66",x"C0",x"C0",x"C0",x"66",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"CC",x"C6",x"C6",x"C6",x"CC",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"3E",x"60",x"C0",x"DE",x"C6",x"66",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"18",x"18",x"18",x"18",x"18",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1E",x"06",x"06",x"06",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"CC",x"D8",x"F0",x"F8",x"DC",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"C6",x"C6",x"C6",x"FC",x"C0",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"DE",x"CC",x"7A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FC",x"C6",x"C6",x"CE",x"F8",x"DC",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"CC",x"C0",x"7C",x"06",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"EE",x"7C",x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"C6",x"C6",x"D6",x"FE",x"FE",x"EE",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"0E",x"1C",x"38",x"70",x"E0",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"0E",x"08",x"08",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"65",x"79",x"65",x"65",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E4",x"96",x"96",x"97",x"96",x"E6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"00",x"59",x"59",x"59",x"59",x"D9",x"4E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"70",x"70",x"3C",x"0C",x"78",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"EE",x"28",x"28",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"0E",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"28",x"28",x"EE",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"70",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"3E",x"3C",x"38",x"30",x"00",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"70",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"FF",x"81",x"81",x"81",x"FF",x"81",x"81",
															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"81",x"FF",x"81",x"81",x"81",x"FF",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"81",x"FF",x"81",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"81",x"FF",x"81",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"C6",x"81",x"FF",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"81",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"38",x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",
															x"6C",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"81",x"81",x"C6",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"FF",x"81",x"81",x"83",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"FF",x"81",x"81",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"81",x"81",x"81",x"FF",x"81",x"81",x"BF",x"5F",x"5F",x"5F",x"00",x"5F",x"51",x"55",x"FF",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"51",x"5F",x"00",x"5F",x"5F",x"5F",x"5F",x"BF",x"7F",x"7F",x"7F",x"7F",x"72",x"7F",x"7F",x"FF",x"FF",x"FE",x"FE",x"FE",x"00",x"FE",x"26",x"26",x"FF",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"22",x"FE",x"00",x"FE",x"FE",x"FE",x"FE",x"FF",x"FE",x"FE",x"FE",x"FE",x"4A",x"FE",x"FE",x"FF",
															x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"05",x"0F",x"0B",x"1B",x"13",x"13",x"13",x"13",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",x"13",x"13",x"13",x"13",x"1B",x"0B",x"0F",x"05",x"07",x"00",x"0F",x"1F",x"1F",x"1F",x"1F",x"1F",x"05",x"0F",x"0B",x"1B",x"13",x"13",x"13",x"13",x"1F",x"1F",x"1F",x"1F",x"1F",x"0F",x"00",x"07",x"13",x"13",x"13",x"13",x"1B",x"0B",x"0F",x"05",x"E0",x"00",x"F1",x"FB",x"FB",x"FB",x"FB",x"FB",x"A0",x"F1",x"D1",x"DB",x"CA",x"CA",x"CA",x"CA",x"FB",x"FB",x"FB",x"FB",x"FB",x"F1",x"00",x"E0",x"CA",x"CA",x"CA",x"CA",x"DB",x"D1",x"F1",x"A0",x"E0",x"00",x"F1",x"FB",x"FB",x"FB",x"FB",x"FB",x"A0",x"F1",x"D1",x"DB",x"CA",x"CA",x"CA",x"CA",x"FB",x"FB",x"FB",x"FB",x"FB",x"F1",x"00",x"E0",x"CA",x"CA",x"CA",x"CA",x"DB",x"D1",x"F0",x"A0",
															x"FC",x"00",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"B4",x"FE",x"7A",x"7B",x"79",x"79",x"79",x"79",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"00",x"FC",x"79",x"79",x"79",x"79",x"7B",x"7A",x"FE",x"B4",x"FC",x"00",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"B4",x"FE",x"7A",x"7B",x"79",x"79",x"79",x"79",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"00",x"FC",x"79",x"79",x"79",x"79",x"7B",x"7A",x"FE",x"B4",x"00",x"00",x"1F",x"10",x"10",x"1F",x"00",x"00",x"7F",x"BF",x"FF",x"B2",x"B1",x"FF",x"BF",x"7F",x"00",x"00",x"F8",x"08",x"08",x"F8",x"00",x"00",x"FE",x"FD",x"FF",x"CD",x"6D",x"FF",x"FD",x"FE",x"00",x"01",x"02",x"02",x"F1",x"08",x"04",x"03",x"FF",x"FF",x"AE",x"FE",x"FF",x"0F",x"07",x"03",x"00",x"80",x"40",x"40",x"8F",x"10",x"20",x"C0",x"FF",x"FF",x"75",x"7F",x"FF",x"F0",x"E0",x"C0",
															x"03",x"04",x"08",x"F1",x"02",x"02",x"01",x"00",x"03",x"07",x"0F",x"FF",x"FE",x"AE",x"FF",x"FF",x"C0",x"20",x"10",x"8F",x"40",x"40",x"80",x"00",x"C0",x"E0",x"F0",x"FF",x"7F",x"75",x"FF",x"FF",x"FF",x"FF",x"C3",x"81",x"81",x"C3",x"FF",x"FF",x"FF",x"00",x"C3",x"81",x"81",x"C3",x"FF",x"00",x"FF",x"99",x"00",x"00",x"00",x"81",x"81",x"81",x"81",x"66",x"7E",x"7E",x"7E",x"FF",x"FF",x"7E",x"00",x"00",x"00",x"00",x"60",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6C",x"6C",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"66",x"66",x"66",x"66",x"66",x"66",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"83",x"D1",x"E1",x"D1",x"02",x"84",x"F0",x"CE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"C1",x"8B",x"87",x"8B",x"40",x"21",x"0F",x"D3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"0F",x"1E",x"3F",x"7F",x"FF",x"FF",x"FF",x"1F",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"F8",x"F0",x"78",x"FC",x"FE",x"FF",x"FF",x"FF",x"F8",x"F8",x"FC",x"FE",x"FF",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"81",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"81",x"81",x"BD",x"7E",x"FF",x"E7",x"FF",x"FF",x"FF",x"81",x"BD",x"7E",x"A5",x"DB",x"E7",x"FF",x"FF",
															x"01",x"07",x"1F",x"3F",x"7F",x"FF",x"FF",x"DD",x"00",x"05",x"19",x"33",x"63",x"C7",x"C7",x"C4",x"89",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"80",x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"80",x"E0",x"F8",x"FC",x"FE",x"FF",x"FF",x"3B",x"00",x"A0",x"98",x"CC",x"C6",x"E3",x"E3",x"23",x"11",x"00",x"00",x"00",x"00",x"40",x"80",x"00",x"01",x"00",x"00",x"00",x"00",x"40",x"80",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"01",x"03",x"00",x"00",x"03",x"19",x"00",x"00",x"01",x"03",x"03",x"07",x"04",x"1C",x"3F",x"7F",x"00",x"00",x"7C",x"02",x"01",x"00",x"00",x"00",x"7F",x"FF",x"FF",x"7F",x"7F",x"1F",x"03",x"00",
															x"00",x"00",x"01",x"01",x"03",x"07",x"07",x"0F",x"00",x"00",x"01",x"01",x"03",x"07",x"07",x"0F",x"0F",x"07",x"0F",x"07",x"01",x"10",x"20",x"00",x"FF",x"FF",x"3F",x"3F",x"7F",x"FE",x"FC",x"30",x"F8",x"FE",x"7F",x"1F",x"0F",x"19",x"30",x"70",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"73",x"27",x"0F",x"1F",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FE",x"FD",x"F8",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"EF",x"CF",x"9F",x"1F",x"0F",x"2D",x"50",x"40",x"EF",x"CF",x"9F",x"1F",x"0F",x"7F",x"FF",x"FF",x"00",x"00",x"00",x"00",x"E0",x"FE",x"FF",x"F3",x"00",x"00",x"00",x"F0",x"FE",x"FF",x"FF",x"FF",x"FB",x"FB",x"FB",x"FB",x"FB",x"F3",x"F7",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"CF",x"9F",x"3F",x"3F",x"3F",x"0F",x"03",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"F0",x"FC",x"F0",x"F0",x"98",x"08",x"00",x"FF",x"FF",x"FF",x"F0",x"F0",x"F8",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",x"F8",x"F8",x"F0",x"F0",x"F8",x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"1F",x"1F",x"0F",x"07",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"0F",x"07",x"00",x"00",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",x"F0",x"F8",x"00",x"80",x"C0",x"E0",x"F0",x"F0",x"F0",x"FC",x"F9",x"FF",x"FF",x"FF",x"FF",x"0E",x"02",x"14",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",x"1F",x"3F",
															x"80",x"A0",x"20",x"20",x"A0",x"80",x"00",x"00",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"C0",x"80",x"01",x"05",x"04",x"04",x"05",x"01",x"00",x"00",x"03",x"07",x"07",x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"03",x"07",x"0F",x"0F",x"0F",x"0F",x"00",x"01",x"03",x"07",x"0F",x"0F",x"0F",x"3F",x"9F",x"FF",x"FF",x"FF",x"FF",x"70",x"40",x"28",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"F8",x"FC",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"1F",x"1F",x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"F8",x"F8",x"F0",x"E0",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"F0",x"E0",x"00",x"00",x"00",
															x"00",x"00",x"00",x"00",x"07",x"7F",x"FF",x"CF",x"00",x"00",x"00",x"0F",x"7F",x"FF",x"FF",x"FF",x"DF",x"DF",x"DF",x"DF",x"DF",x"CF",x"EF",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F3",x"F9",x"FC",x"FC",x"FC",x"F0",x"C0",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"0F",x"3F",x"0F",x"0F",x"19",x"10",x"00",x"FF",x"FF",x"FF",x"0F",x"0F",x"1F",x"1F",x"1F",x"1F",x"7F",x"FE",x"F8",x"F0",x"98",x"0C",x"0E",x"1F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"CE",x"E4",x"F0",x"F8",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"7F",x"BF",x"1F",x"6F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F7",x"F3",x"F9",x"F8",x"F0",x"B4",x"0A",x"02",x"F7",x"F3",x"F9",x"F8",x"F0",x"FE",x"FF",x"FF",
															x"80",x"C0",x"00",x"00",x"C0",x"98",x"00",x"00",x"80",x"C0",x"C0",x"E0",x"20",x"38",x"FC",x"FE",x"00",x"00",x"3E",x"40",x"80",x"00",x"00",x"00",x"FE",x"FF",x"FF",x"FE",x"FC",x"F8",x"C0",x"00",x"00",x"00",x"80",x"80",x"C0",x"E0",x"E0",x"F0",x"00",x"00",x"80",x"80",x"C0",x"E0",x"E0",x"F0",x"F0",x"E0",x"F0",x"E0",x"80",x"08",x"04",x"00",x"FF",x"FF",x"FC",x"FC",x"FE",x"7E",x"3F",x"0C",x"00",x"00",x"01",x"03",x"03",x"03",x"07",x"07",x"00",x"01",x"03",x"07",x"07",x"07",x"0F",x"0F",x"07",x"03",x"03",x"03",x"03",x"03",x"03",x"01",x"0F",x"0F",x"07",x"07",x"07",x"03",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"01",x"01",x"01",x"00",x"00",x"03",x"07",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"1C",x"3B",x"00",x"00",x"00",x"00",x"01",x"03",x"3F",x"7F",
															x"7E",x"FE",x"FF",x"FF",x"FF",x"FF",x"FD",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"F9",x"F3",x"F7",x"F6",x"EE",x"FD",x"FC",x"F8",x"E1",x"F3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D3",x"CB",x"C3",x"E1",x"F9",x"39",x"42",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"07",x"0F",x"19",x"30",x"63",x"72",x"70",x"01",x"07",x"0F",x"1F",x"3F",x"FC",x"FC",x"FF",x"FF",x"00",x"1F",x"20",x"C0",x"C0",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"AB",x"C1",x"81",x"91",x"82",x"FC",x"E0",x"CE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E5",x"DA",x"F0",x"E0",x"C0",x"00",x"00",x"00",x"FF",x"FF",x"F0",x"E0",x"C0",x"80",x"80",x"00",x"F0",x"F8",x"CC",x"86",x"62",x"26",x"06",x"C0",x"F0",x"F8",x"FC",x"FE",x"9F",x"9F",x"FF",x"FF",
															x"00",x"FC",x"06",x"03",x"01",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D5",x"83",x"81",x"89",x"41",x"3F",x"07",x"D3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"6F",x"DB",x"0F",x"07",x"03",x"00",x"00",x"00",x"FF",x"FF",x"0F",x"07",x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"DC",x"00",x"00",x"00",x"00",x"80",x"C0",x"FC",x"FE",x"7E",x"7F",x"7F",x"FF",x"FF",x"FF",x"BF",x"9F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BF",x"9F",x"CF",x"EF",x"6F",x"77",x"BF",x"3F",x"1F",x"87",x"CF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CB",x"D3",x"C3",x"87",x"9F",x"9C",x"42",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"80",x"C0",x"C0",x"C0",x"E0",x"E0",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"F0",x"F0",
															x"E0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"80",x"F0",x"F0",x"E0",x"E0",x"E0",x"C0",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",x"80",x"40",x"20",x"80",x"80",x"80",x"00",x"00",x"C0",x"E0",x"F0",x"00",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"00",x"00",x"01",x"03",x"07",x"07",x"07",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"01",x"01",x"03",x"01",x"00",x"00",x"00",x"01",x"03",x"03",x"01",x"01",x"07",x"03",x"04",x"00",x"00",x"00",x"03",x"03",x"07",x"1F",x"3F",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"01",x"03",x"03",x"0F",x"0E",x"3E",x"7F",x"FF",x"FF",x"EF",x"F7",x"F8",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"1F",x"1F",x"7F",x"FF",x"FE",x"FF",x"FF",x"FF",x"1F",x"7F",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FC",x"F8",x"80",x"00",x"00",x"FF",x"FF",x"FF",x"FC",x"F8",x"F8",x"00",x"00",x"30",x"7F",x"7F",x"3F",x"87",x"F0",x"FF",x"FF",x"CF",x"88",x"DD",x"C8",x"F8",x"FF",x"FF",x"FF",x"E5",x"DA",x"C0",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"C0",x"00",x"00",x"00",x"00",x"00",x"06",x"FF",x"FF",x"FE",x"F1",x"07",x"FF",x"FF",x"F9",x"88",x"DD",x"89",x"0F",x"FF",x"FF",x"FF",x"00",x"01",x"02",x"07",x"00",x"00",x"20",x"FF",x"03",x"07",x"0F",x"07",x"87",x"C3",x"E0",x"FF",x"7F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"B8",x"78",x"78",x"B0",x"78",x"FC",x"FE",x"FC",x"F8",x"F8",x"F8",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"9C",x"42",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"00",x"00",x"20",x"40",x"8A",x"1E",x"7E",x"BE",x"C0",x"F0",x"FC",x"FC",x"FE",x"FE",x"FE",x"FE",x"DF",x"FF",x"FE",x"FC",x"F0",x"E0",x"80",x"00",x"FF",x"FF",x"FE",x"FC",x"F0",x"E0",x"80",x"00",x"00",x"00",x"04",x"02",x"51",x"78",x"7E",x"FD",x"03",x"0F",x"3F",x"3F",x"7F",x"7F",x"7E",x"FF",x"FB",x"FF",x"7F",x"3F",x"0F",x"07",x"01",x"00",x"FF",x"FF",x"7F",x"3F",x"0F",x"07",x"01",x"00",x"00",x"80",x"40",x"E0",x"00",x"00",x"04",x"FF",x"C0",x"E0",x"F0",x"E0",x"E1",x"C3",x"07",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1D",x"1E",x"1E",x"0D",x"1E",x"3F",x"7F",x"3F",x"1F",x"1F",x"1F",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"39",x"42",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"6F",x"DB",x"03",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"00",x"00",x"00",x"00",x"80",x"C0",x"C0",x"F0",x"70",x"7C",x"7E",x"FF",x"FF",x"F7",x"EF",x"1F",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"1E",x"01",x"00",x"00",x"FF",x"FF",x"FF",x"3F",x"1F",x"1F",x"00",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"00",x"00",x"80",x"C0",x"E0",x"E0",x"E0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",x"80",x"80",x"C0",x"80",x"00",x"00",x"00",x"80",x"C0",x"C0",x"80",x"80",x"E0",x"C0",x"20",x"00",x"00",x"00",x"C0",x"C0",x"E0",x"F8",x"FC",x"FC",x"00",x"00",
															x"1F",x"06",x"06",x"06",x"06",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"39",x"65",x"65",x"65",x"65",x"65",x"39",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"B0",x"B0",x"B6",x"E6",x"80",x"80",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"01",x"07",x"00",x"00",x"00",x"00",x"03",x"07",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"7F",x"7F",x"FF",x"7F",x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"7F",x"00",x"00",x"00",x"80",x"00",x"00",x"00",x"A0",x"00",x"00",x"00",x"C0",x"E0",x"F0",x"F0",x"F8",x"E0",x"F0",x"E0",x"DD",x"FA",x"EB",x"80",x"00",x"FC",x"F8",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"00",x"00",x"00",x"03",x"06",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"03",x"07",x"0F",x"1F",x"0B",x"07",x"03",x"5D",x"AF",x"53",x"00",x"00",x"3F",x"1F",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"80",x"00",x"00",x"60",x"F0",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"E0",x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FF",x"FF",x"7E",x"FC",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"21",x"3F",x"36",x"36",x"7E",x"7F",x"7F",x"7F",x"3F",x"3F",x"3F",x"1F",x"1F",x"0F",x"07",x"03",x"00",x"00",x"3F",x"1F",x"1F",x"0F",x"07",x"03",x"00",x"00",x"3E",x"1E",x"1E",x"0E",x"0F",x"1F",x"9F",x"9F",x"3F",x"1F",x"DF",x"CF",x"CF",x"9F",x"DF",x"FF",x"DF",x"FF",x"FF",x"FF",x"FF",x"DF",x"E7",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"0F",
															x"20",x"0F",x"30",x"40",x"98",x"3E",x"1F",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"81",x"36",x"2E",x"AF",x"AE",x"D1",x"EF",x"87",x"FF",x"F9",x"F0",x"F0",x"B1",x"DF",x"EF",x"87",x"02",x"F8",x"06",x"01",x"0C",x"3E",x"FC",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"36",x"3E",x"7A",x"B6",x"CD",x"FB",x"F0",x"FF",x"CF",x"87",x"87",x"CE",x"FD",x"FB",x"F0",x"3E",x"3C",x"3C",x"38",x"F8",x"7C",x"7E",x"78",x"FE",x"FC",x"FC",x"F8",x"FB",x"FD",x"FE",x"FF",x"F8",x"7F",x"7F",x"FE",x"FF",x"FF",x"F3",x"81",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"00",x"00",x"00",x"10",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"78",x"FC",x"FC",x"FC",x"FC",x"06",x"0E",x"7E",x"FE",x"FE",x"FC",x"F8",x"F0",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"F8",x"F0",
															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"08",x"01",x"13",x"01",x"00",x"00",x"01",x"0F",x"1F",x"1F",x"3B",x"33",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"6C",x"FD",x"FF",x"FF",x"00",x"43",x"7F",x"7F",x"7F",x"3F",x"1F",x"07",x"FF",x"7F",x"7F",x"7F",x"7F",x"3F",x"1F",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"10",x"38",x"BF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"7E",x"1E",x"1E",x"0E",x"0F",x"1E",x"1E",x"3E",x"FF",x"7F",x"1F",x"0F",x"0F",x"9F",x"9F",x"BF",x"7F",x"7F",x"BF",x"FF",x"FF",x"FF",x"E7",x"C0",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"CF",
															x"00",x"00",x"10",x"FD",x"FA",x"EB",x"80",x"00",x"00",x"00",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"20",x"1F",x"60",x"8E",x"3F",x"7F",x"7F",x"7C",x"FF",x"FF",x"FF",x"F1",x"C4",x"EE",x"C4",x"83",x"39",x"36",x"2E",x"AF",x"AE",x"D1",x"EF",x"87",x"C7",x"F9",x"F0",x"F0",x"B1",x"DF",x"EF",x"87",x"00",x"00",x"04",x"5F",x"AF",x"53",x"00",x"00",x"00",x"00",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"02",x"FC",x"03",x"38",x"FE",x"FF",x"FF",x"1E",x"FF",x"FF",x"FF",x"C7",x"45",x"EE",x"44",x"E1",x"C0",x"36",x"3E",x"7A",x"B6",x"CD",x"FB",x"F0",x"FF",x"CF",x"87",x"87",x"CE",x"FD",x"FB",x"F0",x"00",x"00",x"00",x"00",x"00",x"0E",x"08",x"08",x"00",x"00",x"00",x"00",x"00",x"01",x"07",x"0F",x"1F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"3F",x"3E",x"3C",x"B8",x"78",x"78",x"7E",x"7E",x"FF",x"FF",x"FD",x"F8",x"FF",x"FF",x"FE",x"FF",x"FD",x"79",x"7B",x"FF",x"FF",x"FF",x"F3",x"80",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"F0",x"10",x"84",x"E0",x"C0",x"80",x"80",x"00",x"00",x"FC",x"FE",x"EC",x"E0",x"C0",x"C0",x"80",x"80",x"00",x"48",x"20",x"00",x"00",x"04",x"0E",x"FE",x"70",x"FC",x"FC",x"FC",x"FC",x"FC",x"FE",x"FE",x"FE",x"FC",x"FC",x"F8",x"F0",x"E0",x"80",x"00",x"FE",x"FC",x"FC",x"F8",x"F0",x"E0",x"80",x"00",x"0F",x"06",x"06",x"06",x"06",x"06",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"60",x"60",x"66",x"66",x"60",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
	
	constant MARIO_BROS_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"00", x"03", x"03", x"0F", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"1F", x"00", x"00", x"00", x"80", x"E0", x"F0", x"F0", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F8", x"04", x"1E", x"00", x"00", x"01", x"03", x"0F", x"1F", x"3F", x"1F", x"0F", x"07", x"20", x"70", x"70", x"20", x"48", x"9C", x"08", x"00", x"F0", x"FC", x"FC", x"F8", x"F8", x"FC", x"F8", x"E0", x"10", x"10", x"32", x"26", x"0F", x"07", x"2F", x"3F", x"1F", x"08", x"00", x"00", x"00", x"04", x"0F", x"0F", x"07", x"00", x"00", x"00", x"F8", x"F8", x"F8", x"F8", x"FE", x"7E", x"06", x"0C", x"7C", x"F8", x"F8", x"F8", x"FC", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"1F", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", 
															x"04", x"08", x"3D", x"00", x"00", x"07", x"0F", x"1F", x"3F", x"7F", x"3F", x"1F", x"0F", x"01", x"C2", x"C2", x"90", x"90", x"38", x"10", x"00", x"E0", x"F0", x"F8", x"F0", x"F0", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"3F", x"7B", x"1F", x"1F", x"0F", x"0F", x"07", x"0F", x"C6", x"07", x"1F", x"1F", x"0F", x"0F", x"00", x"00", x"F0", x"E0", x"E0", x"F4", x"FE", x"7A", x"00", x"00", x"0C", x"1C", x"FC", x"F8", x"F8", x"78", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"0F", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"1F", x"00", x"00", x"00", x"80", x"E0", x"F0", x"F0", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F8", x"04", x"1E", x"00", x"00", x"03", x"07", x"0F", x"0F", x"3F", x"1F", x"0F", x"07", x"00", x"01", x"01", x"33", x"48", x"9C", x"08", x"00", x"E0", x"F0", x"F8", x"F8", x"F8", x"FC", x"F8", x"E0", x"80", x"00", x"00", x"C0", 
															x"0D", x"0D", x"0B", x"07", x"07", x"0F", x"00", x"00", x"3F", x"3F", x"0F", x"07", x"00", x"00", x"00", x"00", x"F8", x"30", x"10", x"30", x"F0", x"E0", x"E0", x"E0", x"80", x"C0", x"F0", x"F0", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"0F", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"1F", x"00", x"00", x"00", x"80", x"E0", x"F0", x"F0", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F8", x"04", x"1E", x"00", x"00", x"07", x"0F", x"3F", x"7F", x"3F", x"1F", x"0F", x"07", x"04", x"08", x"08", x"08", x"88", x"1C", x"08", x"00", x"F0", x"FC", x"FE", x"FE", x"F8", x"FC", x"F8", x"E0", x"60", x"60", x"C0", x"81", x"34", x"1F", x"1F", x"1F", x"3F", x"3C", x"38", x"78", x"DF", x"FF", x"5F", x"1F", x"3F", x"3C", x"00", x"00", x"F4", x"F0", x"F0", x"F8", x"FC", x"3C", x"1C", x"1E", x"F3", x"F7", x"F2", x"F8", x"FC", x"3C", x"00", x"00", 
															x"00", x"00", x"00", x"10", x"18", x"3B", x"38", x"38", x"00", x"1C", x"1E", x"0E", x"04", x"00", x"00", x"07", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"3C", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FE", x"31", x"3F", x"1C", x"1E", x"0F", x"0F", x"4F", x"4F", x"0F", x"07", x"03", x"03", x"06", x"0C", x"09", x"0F", x"12", x"A7", x"02", x"00", x"FC", x"FE", x"FC", x"F0", x"FE", x"FF", x"FE", x"F8", x"60", x"C0", x"83", x"87", x"7E", x"7F", x"7F", x"07", x"00", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"07", x"00", x"00", x"00", x"00", x"F0", x"F8", x"FC", x"FE", x"F2", x"60", x"00", x"00", x"D2", x"F0", x"E0", x"F0", x"F0", x"60", x"00", x"00", x"03", x"0F", x"00", x"02", x"04", x"1E", x"00", x"7F", x"00", x"00", x"03", x"1F", x"3F", x"1F", x"0F", x"04", x"E0", x"F0", x"F0", x"48", x"48", x"9C", x"08", x"FE", x"00", x"00", x"F0", x"F8", x"F8", x"FC", x"F8", x"40", 
															x"FF", x"37", x"1F", x"1F", x"3F", x"3F", x"3C", x"78", x"08", x"DF", x"DF", x"1F", x"3F", x"3F", x"3C", x"00", x"FF", x"78", x"F8", x"F8", x"FC", x"FC", x"3C", x"1E", x"80", x"E7", x"FB", x"F8", x"FC", x"FC", x"3C", x"00", x"00", x"00", x"00", x"03", x"0F", x"02", x"04", x"1E", x"00", x"00", x"00", x"00", x"00", x"1F", x"3F", x"1F", x"00", x"00", x"00", x"E0", x"F0", x"78", x"24", x"46", x"00", x"00", x"00", x"00", x"00", x"F8", x"FC", x"FE", x"00", x"7F", x"FF", x"37", x"1F", x"3F", x"3F", x"78", x"0F", x"0C", x"08", x"DF", x"DF", x"3F", x"3F", x"00", x"08", x"FC", x"FF", x"7C", x"F8", x"FC", x"FC", x"1E", x"F8", x"60", x"C0", x"C3", x"FF", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"1C", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FE", 
															x"01", x"07", x"00", x"00", x"03", x"07", x"7F", x"7F", x"0F", x"07", x"03", x"31", x"78", x"74", x"09", x"1B", x"12", x"E7", x"C2", x"00", x"FC", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"F8", x"30", x"40", x"80", x"80", x"3D", x"1F", x"0F", x"5F", x"5F", x"7F", x"3C", x"10", x"3F", x"1F", x"0F", x"1F", x"1F", x"0F", x"04", x"00", x"F7", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"90", x"DF", x"F7", x"E4", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"1C", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FE", x"01", x"07", x"00", x"00", x"03", x"07", x"7F", x"7F", x"0F", x"07", x"03", x"31", x"78", x"74", x"09", x"1B", x"12", x"E7", x"C2", x"00", x"FC", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"F8", x"30", x"40", x"80", x"80", 
															x"3D", x"1F", x"0F", x"5F", x"5F", x"7F", x"3C", x"10", x"3F", x"1F", x"0F", x"1F", x"1F", x"0F", x"04", x"01", x"F7", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"90", x"DF", x"FF", x"E4", x"C0", x"10", x"40", x"00", x"00", x"02", x"17", x"0F", x"01", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"06", x"07", x"0F", x"3F", x"00", x"00", x"00", x"80", x"C0", x"E0", x"E0", x"90", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"08", x"3C", x"00", x"00", x"3F", x"3F", x"3F", x"1F", x"7F", x"3D", x"01", x"3F", x"C8", x"D0", x"D1", x"59", x"10", x"38", x"10", x"7C", x"FC", x"FC", x"F0", x"F8", x"F0", x"F8", x"F0", x"83", x"83", x"83", x"82", x"88", x"16", x"0F", x"0F", x"07", x"03", x"00", x"00", x"00", x"1F", x"0F", x"0F", x"07", x"03", x"00", x"00", x"00", x"F8", x"FE", x"FF", x"FF", x"FF", x"E2", x"60", x"00", x"D8", x"FC", x"FC", x"FC", x"F8", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"07", x"0F", x"10", x"12", x"02", x"00", x"00", x"00", x"01", x"00", x"1F", x"5F", x"DF", x"00", x"60", x"F0", x"F0", x"F0", x"10", x"90", x"80", x"00", x"60", x"90", x"00", x"00", x"F0", x"F4", x"F7", x"28", x"3C", x"37", x"30", x"10", x"18", x"3C", x"3F", x"DF", x"4F", x"0F", x"0F", x"0C", x"0C", x"3B", x"3C", x"28", x"7C", x"D8", x"18", x"10", x"30", x"7C", x"FC", x"F7", x"E0", x"E0", x"E0", x"60", x"60", x"BC", x"7C", x"FB", x"FF", x"FF", x"77", x"33", x"00", x"00", x"00", x"3F", x"1F", x"1F", x"07", x"03", x"00", x"00", x"00", x"BF", x"FF", x"FF", x"EE", x"CC", x"00", x"00", x"00", x"FC", x"F8", x"F8", x"E0", x"C0", x"00", x"00", x"00", x"00", x"07", x"05", x"01", x"03", x"06", x"04", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"04", x"04", x"07", x"01", x"05", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"07", x"05", x"05", x"07", x"05", x"05", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"27", x"25", x"25", x"25", x"25", x"25", x"27", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"27", x"24", x"24", x"27", x"25", x"25", x"27", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"75", x"55", x"15", x"35", x"67", x"41", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"77", x"55", x"11", x"33", x"16", x"54", x"77", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"77", x"55", x"55", x"55", x"55", x"55", x"77", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"38", x"54", x"FE", x"54", x"38", x"10", x"00", x"00", x"28", x"6C", x"00", x"6C", x"28", x"00", x"00", x"38", x"7C", x"C6", x"C6", x"C6", x"7C", x"38", x"00", x"38", x"6C", x"FE", x"BA", x"FE", x"6C", x"38", x"00", 
															x"10", x"54", x"28", x"C6", x"28", x"54", x"10", x"00", x"00", x"10", x"38", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"01", x"10", x"00", x"00", x"01", x"23", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"10", x"00", x"00", x"00", x"88", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"01", x"00", x"00", x"10", x"01", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"14", x"3E", x"55", x"54", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"15", x"55", x"3E", x"14", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"18", x"18", x"30", x"00", x"00", x"00", x"00", x"00", x"04", x"46", x"4E", x"FE", x"FE", x"EC", x"5C", x"1C", x"26", x"5B", x"A5", x"DB", x"66", x"3C", x"00", x"F8", x"E4", x"DA", x"A5", x"DB", x"66", x"7E", x"E7", x"1C", x"0C", x"0C", x"18", x"00", x"00", x"00", x"00", x"00", x"22", x"63", x"E7", x"FF", x"4F", x"0E", x"1C", x"1C", x"26", x"5B", x"A5", x"DB", x"7C", x"00", x"00", x"F8", x"E4", x"DA", x"A5", x"DB", x"7E", x"47", x"E0", x"1C", x"0C", x"0C", x"18", x"00", x"00", x"00", x"00", x"00", x"02", x"23", x"67", x"7F", x"7F", x"26", x"0E", x"1C", x"26", x"5B", x"A5", x"DB", x"3E", x"00", x"00", x"78", x"64", x"DA", x"A5", x"DB", x"7E", x"E2", x"07", 
															x"18", x"30", x"30", x"38", x"10", x"00", x"00", x"00", x"04", x"06", x"47", x"47", x"6D", x"7C", x"3E", x"1C", x"20", x"70", x"A8", x"DC", x"AA", x"77", x"2B", x"1E", x"EC", x"F8", x"A9", x"DF", x"AA", x"77", x"2A", x"18", x"18", x"30", x"30", x"38", x"10", x"00", x"00", x"00", x"26", x"47", x"45", x"40", x"68", x"78", x"3E", x"1C", x"20", x"70", x"A8", x"DC", x"AA", x"77", x"2B", x"1E", x"F0", x"F8", x"AB", x"DE", x"AA", x"77", x"2A", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6A", x"DB", x"A5", x"DB", x"66", x"3C", x"A2", x"D6", x"FE", x"DB", x"A5", x"DA", x"64", x"38", x"00", x"00", x"5C", x"DB", x"A5", x"DB", x"62", x"3C", x"00", x"00", x"5C", x"DB", x"A5", x"DA", x"60", x"38", x"00", x"00", x"6E", x"DB", x"A5", x"DB", x"62", x"3C", x"00", x"00", x"6E", x"DB", x"A5", x"DA", x"60", x"38", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"08", x"1D", x"12", x"20", x"01", x"00", x"00", x"00", x"07", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"A6", x"D0", x"98", x"04", x"00", x"00", x"00", x"F0", x"50", x"00", x"00", x"00", x"00", x"00", x"00", x"33", x"71", x"28", x"3F", x"71", x"40", x"80", x"01", x"0F", x"0F", x"17", x"00", x"00", x"00", x"00", x"00", x"E4", x"06", x"6D", x"68", x"96", x"8D", x"80", x"00", x"F8", x"F8", x"90", x"90", x"08", x"00", x"00", x"00", x"00", x"26", x"56", x"54", x"F4", x"F6", x"62", x"3A", x"30", x"60", x"D0", x"D0", x"F0", x"F0", x"62", x"3A", x"00", x"C8", x"D4", x"5A", x"5F", x"CF", x"86", x"9C", x"00", x"0C", x"16", x"1B", x"1F", x"0F", x"86", x"9C", x"FF", x"56", x"7E", x"7E", x"3C", x"A5", x"A5", x"A5", x"FB", x"54", x"7E", x"7E", x"BD", x"A5", x"A5", x"A5", x"00", x"06", x"16", x"24", x"2C", x"7E", x"72", x"1A", x"00", x"18", x"30", x"60", x"68", x"78", x"72", x"1A", 
															x"08", x"C6", x"E6", x"73", x"5B", x"DF", x"8E", x"9C", x"0C", x"04", x"27", x"33", x"1B", x"1F", x"8E", x"9C", x"FF", x"56", x"7E", x"7E", x"3C", x"95", x"5A", x"50", x"FB", x"54", x"7E", x"7F", x"BC", x"95", x"5A", x"50", x"06", x"36", x"24", x"6C", x"7E", x"7A", x"32", x"1F", x"38", x"70", x"60", x"68", x"78", x"7A", x"32", x"1F", x"D8", x"CC", x"64", x"76", x"DE", x"8C", x"98", x"F0", x"1C", x"0E", x"26", x"36", x"1E", x"8C", x"98", x"B0", x"D7", x"7E", x"7E", x"7E", x"95", x"95", x"49", x"02", x"D5", x"7E", x"7E", x"FF", x"95", x"95", x"49", x"02", x"14", x"34", x"34", x"36", x"3E", x"3E", x"1C", x"08", x"14", x"36", x"36", x"36", x"3E", x"3E", x"1C", x"08", x"0C", x"1C", x"34", x"3C", x"7D", x"41", x"41", x"22", x"18", x"3C", x"34", x"3E", x"3D", x"41", x"41", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"18", x"05", x"03", x"05", x"07", x"07", x"0C", x"1F", x"07", x"1A", x"0F", x"07", x"07", x"06", x"00", x"00", x"0C", x"D0", x"E0", x"D0", x"F0", x"70", x"38", x"7C", x"70", x"2C", x"78", x"70", x"70", x"B0", x"14", x"55", x"BD", x"3C", x"3C", x"18", x"C3", x"00", x"2A", x"2A", x"3C", x"00", x"7E", x"5A", x"C3", x"00", 
															x"00", x"00", x"18", x"05", x"03", x"05", x"07", x"07", x"00", x"30", x"64", x"6A", x"7B", x"3F", x"1F", x"06", x"00", x"00", x"0C", x"D0", x"E0", x"D0", x"F0", x"70", x"00", x"0E", x"13", x"2B", x"6F", x"7E", x"7C", x"B0", x"94", x"55", x"3E", x"3C", x"3C", x"D8", x"00", x"03", x"2A", x"2A", x"3C", x"40", x"7C", x"DE", x"02", x"03", x"00", x"00", x"00", x"00", x"03", x"05", x"07", x"07", x"00", x"00", x"00", x"30", x"3B", x"6F", x"7F", x"3E", x"00", x"00", x"00", x"00", x"E0", x"D0", x"F0", x"70", x"00", x"00", x"00", x"06", x"6F", x"7B", x"7F", x"BC", x"14", x"55", x"BF", x"3C", x"3C", x"18", x"03", x"C0", x"EB", x"2A", x"3E", x"00", x"3E", x"7A", x"43", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1F", x"03", x"0F", x"01", x"1F", x"07", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"EC", x"CC", x"44", x"04", x"00", x"00", x"00", x"01", x"13", x"33", x"BB", x"FB", x"FF", x"08", x"08", x"28", x"3A", x"3E", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"28", x"7E", x"FF", x"FF", x"FF", x"FF", x"81", x"FF", x"7E", x"28", x"00", x"28", x"54", x"00", x"7E", x"00", x"00", x"08", x"08", x"28", x"3A", x"36", x"22", x"2A", x"28", x"00", x"00", x"00", x"00", x"08", x"5C", x"7C", x"7E", x"28", x"03", x"AF", x"FF", x"FF", x"81", x"FF", x"7E", x"7E", x"FC", x"78", x"54", x"00", x"7E", x"00", x"00", 
															x"08", x"08", x"28", x"3A", x"36", x"22", x"2A", x"28", x"00", x"00", x"00", x"00", x"08", x"5C", x"7C", x"7E", x"28", x"00", x"28", x"54", x"00", x"00", x"00", x"00", x"7E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"1C", x"36", x"3B", x"33", x"1B", x"0E", x"0C", x"58", x"1C", x"3E", x"37", x"3F", x"1F", x"0E", x"0C", x"58", x"38", x"7C", x"C6", x"AE", x"BB", x"F1", x"60", x"02", x"38", x"7C", x"FE", x"DE", x"FB", x"F1", x"60", x"02", x"34", x"60", x"E0", x"F8", x"DC", x"D6", x"66", x"3C", x"34", x"60", x"E0", x"F8", x"FC", x"EE", x"7E", x"3C", x"40", x"06", x"8F", x"DD", x"75", x"63", x"3E", x"1C", x"40", x"06", x"8F", x"DF", x"7B", x"7F", x"3E", x"1C", x"00", x"00", x"00", x"00", x"07", x"07", x"1F", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", 
															x"3B", x"77", x"02", x"1F", x"0F", x"06", x"CD", x"DD", x"3F", x"7F", x"3F", x"1F", x"0F", x"01", x"C2", x"C2", x"60", x"60", x"C0", x"E0", x"C0", x"E0", x"F0", x"F8", x"F0", x"F0", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"F9", x"7C", x"00", x"00", x"00", x"00", x"07", x"0F", x"C6", x"07", x"1F", x"1F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"18", x"14", x"0C", x"04", x"08", x"00", x"00", x"00", x"18", x"1C", x"0C", x"04", x"08", x"00", x"00", x"00", x"10", x"28", x"10", x"00", x"00", x"00", x"00", x"00", x"10", x"28", x"10", x"00", x"00", x"00", x"00", x"10", x"00", x"54", x"00", x"10", x"00", x"00", x"00", x"10", x"00", x"54", x"00", x"10", x"00", x"00", x"10", x"44", x"10", x"AA", x"10", x"44", x"10", x"00", x"10", x"44", x"10", x"AA", x"10", x"44", x"10", x"00", x"10", x"44", x"00", x"82", x"00", x"44", x"10", x"00", x"10", x"44", x"00", x"82", x"00", x"44", x"10", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"10", x"20", x"20", x"20", x"00", x"00", x"00", x"00", x"18", x"3C", x"1C", x"3C", x"20", x"20", x"20", x"20", x"20", x"20", x"10", x"00", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"00", x"20", x"40", x"80", x"94", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7F", x"FB", x"94", x"94", x"94", x"94", x"48", x"40", x"20", x"00", x"FB", x"FB", x"FB", x"FB", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"38", x"7E", x"FE", x"FE", x"00", x"00", x"00", x"00", x"3C", x"7C", x"FC", x"FF", 
															x"FE", x"FE", x"FE", x"FE", x"7E", x"7E", x"3C", x"00", x"FF", x"FF", x"FF", x"FF", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"08", x"1C", x"1E", x"1E", x"00", x"00", x"00", x"00", x"0C", x"1E", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"18", x"08", x"00", x"1E", x"1E", x"1E", x"1E", x"1E", x"1E", x"0C", x"00", x"30", x"3E", x"1E", x"0E", x"0E", x"06", x"02", x"00", x"CE", x"C2", x"E6", x"EE", x"8E", x"46", x"32", x"0E", x"00", x"00", x"00", x"00", x"02", x"06", x"0E", x"3E", x"00", x"00", x"00", x"02", x"06", x"0A", x"36", x"C6", x"00", x"00", x"3C", x"7E", x"1E", x"0E", x"06", x"02", x"00", x"3C", x"C2", x"86", x"EE", x"EE", x"C6", x"C2", x"00", x"00", x"00", x"00", x"40", x"20", x"30", x"1C", x"00", x"00", x"00", x"C0", x"A0", x"D0", x"CC", x"E2", x"7E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"8E", x"EE", x"E2", x"C4", x"C8", x"B0", x"C0", x"00", 
															x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BE", x"C2", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"0E", x"0E", x"06", x"02", x"02", x"00", x"00", x"E6", x"8E", x"CE", x"26", x"12", x"0E", x"02", x"00", x"00", x"00", x"00", x"3C", x"7E", x"C3", x"81", x"00", x"3C", x"7E", x"FF", x"C3", x"81", x"3C", x"7E", x"FF", x"00", x"81", x"C3", x"FF", x"FF", x"7E", x"3C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"06", x"06", x"0C", x"09", x"19", x"00", x"00", x"00", x"01", x"01", x"03", x"06", x"06", x"80", x"40", x"E0", x"E0", x"A0", x"B0", x"80", x"D0", x"00", x"80", x"00", x"00", x"40", x"40", x"60", x"20", 
															x"08", x"1C", x"3E", x"1F", x"25", x"00", x"02", x"02", x"04", x"02", x"01", x"00", x"0A", x"03", x"01", x"01", x"00", x"70", x"7C", x"F8", x"A0", x"40", x"C0", x"C0", x"70", x"88", x"80", x"00", x"54", x"80", x"00", x"00", x"03", x"06", x"06", x"04", x"0D", x"09", x"19", x"33", x"00", x"01", x"01", x"03", x"02", x"06", x"06", x"0C", x"C0", x"C0", x"E0", x"E0", x"A0", x"B0", x"90", x"48", x"00", x"00", x"00", x"00", x"40", x"40", x"60", x"B0", x"00", x"00", x"30", x"60", x"00", x"00", x"20", x"00", x"00", x"30", x"48", x"80", x"81", x"00", x"00", x"00", x"00", x"00", x"4C", x"00", x"02", x"00", x"00", x"00", x"00", x"0C", x"12", x"02", x"01", x"01", x"00", x"02", x"01", x"03", x"02", x"07", x"06", x"0C", x"19", x"33", x"00", x"00", x"01", x"00", x"01", x"03", x"06", x"0C", x"40", x"C0", x"C0", x"C0", x"E0", x"A0", x"50", x"4C", x"00", x"00", x"00", x"00", x"00", x"40", x"A0", x"B0", 
															x"DB", x"7E", x"5A", x"66", x"34", x"66", x"3C", x"18", x"BD", x"BD", x"BD", x"99", x"5A", x"5A", x"42", x"24", x"18", x"3C", x"00", x"48", x"42", x"E7", x"42", x"40", x"24", x"24", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E3", x"94", x"94", x"E4", x"94", x"94", x"E3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B5", x"B5", x"AD", x"AD", x"AD", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"26", x"29", x"28", x"26", x"21", x"29", x"C6", x"00", x"00", x"20", x"40", x"FE", x"40", x"20", x"00", x"00", x"00", x"20", x"40", x"FE", x"40", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"63", x"94", x"84", x"84", x"84", x"94", x"63", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"29", x"AD", x"AD", x"AB", x"AB", x"AB", x"29", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"34", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"4E", x"2C", x"18", x"00", x"00", x"00", x"00", x"00", x"78", x"30", x"10", x"30", x"78", x"7C", x"78", x"20", x"0E", x"0C", x"08", x"0C", x"06", x"06", x"46", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"EE", x"EE", x"00", x"00", x"EE", x"EE", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"EE", x"00", x"00", x"00", x"00", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"11", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"08", x"04", x"17", x"27", x"55", x"D6", x"72", x"3F", x"08", x"04", x"33", x"61", x"D0", x"D0", x"72", x"3F", x"20", x"40", x"D0", x"C8", x"54", x"D6", x"9E", x"FC", x"20", x"40", x"98", x"0C", x"16", x"16", x"9E", x"BC", x"D7", x"7E", x"D6", x"D6", x"D7", x"24", x"A5", x"A5", x"D5", x"7E", x"C6", x"82", x"01", x"A5", x"A5", x"A5", x"08", x"04", x"27", x"17", x"55", x"F6", x"62", x"3F", x"08", x"24", x"63", x"D1", x"D0", x"F0", x"62", x"3F", x"20", x"48", x"C4", x"CA", x"4B", x"CF", x"9C", x"F0", x"20", x"4C", x"86", x"0B", x"0B", x"0F", x"9C", x"B0", x"D6", x"7E", x"D6", x"D7", x"56", x"95", x"5A", x"50", x"D4", x"7E", x"C6", x"83", x"81", x"95", x"5A", x"50", x"28", x"44", x"57", x"57", x"F5", x"66", x"32", x"1F", x"68", x"C4", x"D3", x"D1", x"F0", x"60", x"32", x"1F", x"24", x"42", x"D2", x"D6", x"5E", x"CC", x"98", x"F0", x"26", x"43", x"93", x"17", x"1E", x"0C", x"98", x"B0", 
															x"D6", x"7E", x"D6", x"D7", x"56", x"95", x"55", x"08", x"D4", x"7E", x"C6", x"83", x"81", x"95", x"55", x"08", x"08", x"24", x"4A", x"10", x"A8", x"AA", x"FE", x"BA", x"08", x"24", x"4A", x"90", x"AA", x"AA", x"FA", x"B8", x"6C", x"5F", x"CF", x"E7", x"7E", x"4E", x"20", x"0E", x"6C", x"5F", x"CF", x"E7", x"70", x"40", x"64", x"60", x"6C", x"DA", x"C7", x"CF", x"EB", x"EB", x"06", x"E0", x"6E", x"FB", x"E7", x"CF", x"0B", x"0B", x"46", x"0C", x"00", x"00", x"00", x"4A", x"91", x"14", x"FE", x"BA", x"00", x"00", x"00", x"4A", x"91", x"55", x"FA", x"B8", x"6C", x"5F", x"CF", x"E7", x"7E", x"4E", x"20", x"0E", x"6C", x"5F", x"CF", x"E7", x"70", x"40", x"64", x"60", x"6C", x"DA", x"C7", x"CF", x"EB", x"EB", x"06", x"E0", x"6E", x"FB", x"E7", x"CF", x"0B", x"0B", x"46", x"0C", x"00", x"00", x"1C", x"7E", x"06", x"25", x"73", x"02", x"00", x"00", x"00", x"00", x"2E", x"FF", x"7F", x"3E", 
															x"00", x"00", x"00", x"00", x"C3", x"00", x"18", x"3C", x"00", x"00", x"00", x"00", x"C3", x"42", x"7E", x"3C", x"03", x"13", x"0A", x"02", x"0E", x"4F", x"3B", x"07", x"00", x"03", x"35", x"75", x"FD", x"BE", x"4E", x"36", x"C0", x"D0", x"A0", x"80", x"E0", x"E4", x"B8", x"C0", x"00", x"C0", x"5C", x"5E", x"7F", x"FB", x"E6", x"D8", x"00", x"00", x"24", x"24", x"00", x"00", x"18", x"3C", x"00", x"00", x"24", x"66", x"42", x"42", x"7E", x"3C", x"03", x"07", x"0A", x"02", x"0E", x"4F", x"3B", x"07", x"38", x"7B", x"E5", x"FD", x"DD", x"3E", x"0E", x"06", x"C0", x"E0", x"90", x"80", x"E0", x"E4", x"B8", x"C0", x"1C", x"DE", x"47", x"7F", x"7A", x"F8", x"E0", x"C0", x"38", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"46", x"C6", x"CF", x"FF", x"F7", x"72", x"3C", x"44", x"6E", x"FF", x"FF", x"FF", x"FF", x"3C", x"00", x"7C", x"7E", x"FF", x"FF", x"E7", x"C3", x"42", x"C3", 
															x"00", x"00", x"22", x"36", x"64", x"8B", x"82", x"C0", x"08", x"08", x"08", x"08", x"1C", x"38", x"55", x"47", x"0E", x"10", x"00", x"00", x"18", x"10", x"18", x"0C", x"06", x"0C", x"19", x"03", x"07", x"0F", x"0E", x"04", x"00", x"00", x"00", x"20", x"58", x"08", x"18", x"30", x"30", x"98", x"D8", x"A0", x"60", x"70", x"E0", x"C0", x"00", x"54", x"60", x"C4", x"15", x"29", x"80", x"00", x"08", x"08", x"00", x"00", x"08", x"1B", x"12", x"40", x"14", x"40", x"00", x"81", x"32", x"40", x"30", x"00", x"0C", x"08", x"00", x"00", x"11", x"3A", x"08", x"00", x"24", x"16", x"00", x"20", x"04", x"02", x"44", x"08", x"00", x"00", x"00", x"00", x"04", x"04", x"68", x"C0", x"92", x"54", x"38", x"FE", x"38", x"54", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"98", x"40", x"02", x"00", x"08", x"00", x"80", x"08", x"80", x"00", x"01", x"02", x"48", x"00", x"00", x"00", x"00", x"20", x"04", x"00", x"01", x"40", x"00", x"10", x"00", x"A0", x"00", x"00", x"00", x"02", x"20", x"00", x"02", x"10", x"00", x"00", x"20", x"02", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"02", x"04", x"26", x"26", x"0E", x"0C", x"1C", x"78", x"F0", x"C0", x"DE", x"DE", x"FE", x"FC", x"FC", x"F8", x"F0", x"C0", x"03", x"0F", x"1D", x"39", x"33", x"63", x"61", x"60", x"03", x"0F", x"1F", x"3F", x"3F", x"7F", x"7F", x"7F", x"C0", x"F0", x"80", x"04", x"01", x"E0", x"F2", x"38", x"C0", x"F0", x"80", x"04", x"01", x"E0", x"F2", x"F8", x"64", x"67", x"63", x"31", x"30", x"18", x"1F", x"0F", x"7B", x"78", x"7C", x"3E", x"3F", x"1F", x"1F", x"0F", x"1C", x"CC", x"CC", x"8C", x"18", x"38", x"F0", x"C0", x"FC", x"3C", x"3C", x"7C", x"F8", x"F8", x"F0", x"C0", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"78", x"C4", x"E4", x"78", x"86", x"86", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"06", x"06", x"06", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"6C", x"6C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"06", x"06", x"06", x"06", x"06", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"60", x"60", x"66", x"66", x"60", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"06", x"06", x"06", x"06", x"06", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"39", x"65", x"65", x"65", x"65", x"65", x"39", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"B0", x"B0", x"B6", x"E6", x"80", x"80", x"00", x"00", x"3C", x"3C", x"00", x"00", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"63", x"63", x"03", x"0E", x"18", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"1F", x"30", x"27", x"2C", x"28", x"28", x"00", x"00", x"00", x"00", x"07", x"0C", x"08", x"08", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"F8", x"0C", x"E4", x"34", x"14", x"14", x"00", x"00", x"00", x"00", x"E0", x"30", x"10", x"10", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"14", x"14", x"14", x"14", x"14", x"14", x"14", x"14", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"28", x"28", x"2C", x"27", x"30", x"1F", x"00", x"00", x"08", x"08", x"0C", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"14", x"14", x"34", x"E4", x"0C", x"F8", x"00", x"00", x"10", x"10", x"30", x"E0", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"80", x"80", x"88", x"88", x"F8", x"FF", x"00", x"00", x"70", x"70", x"7F", x"7F", x"0F", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"8F", x"88", x"88", x"88", x"88", x"88", x"88", x"8F", x"78", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"03", x"01", x"00", x"00", x"00", x"00", x"E0", x"00", x"FC", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"F0", x"78", x"38", x"38", x"38", x"38", x"3C", x"3F", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"88", x"00", x"00", x"00", x"00", x"00", x"00", x"70", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"6F", x"6F", x"6F", x"68", x"60", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"F0", x"F0", x"00", x"00", x"F0", x"F8", x"F8", x"F8", x"78", x"38", x"38", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"C0", x"E0", x"7F", x"3F", x"00", x"00", x"00", x"00", x"3F", x"1F", x"80", x"C0", x"FF", x"FF", x"FF", x"FF", x"88", x"F8", x"FF", x"8F", x"88", x"88", x"88", x"88", x"7F", x"0F", x"08", x"78", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"3C", x"3E", x"3F", x"1F", x"1F", x"0F", x"00", x"00", x"7F", x"7F", x"7F", x"3F", x"3F", x"1F", x"0F", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"88", x"88", x"8F", x"6F", x"6F", x"6F", x"68", x"00", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"F0", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"01", x"01", x"11", x"11", x"1F", x"FF", x"00", x"00", x"0E", x"0E", x"FE", x"FE", x"F0", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F1", x"11", x"11", x"11", x"11", x"11", x"11", x"F1", x"1E", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"C0", x"80", x"00", x"00", x"00", x"00", x"07", x"00", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"0F", x"1E", x"1C", x"1C", x"1C", x"1C", x"3C", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"11", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"FE", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"F6", x"F6", x"F6", x"16", x"06", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"00", x"00", x"0F", x"1F", x"1F", x"1F", x"1E", x"1C", x"1C", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"03", x"07", x"FE", x"FC", x"00", x"00", x"00", x"00", x"FC", x"F8", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"11", x"1F", x"FF", x"F1", x"11", x"11", x"11", x"11", x"FE", x"F0", x"10", x"1E", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7C", x"FC", x"F8", x"F8", x"F0", x"00", x"00", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"F0", x"00", 
															x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"11", x"11", x"F1", x"F6", x"F6", x"F6", x"16", x"00", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"0F", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"00", x"30", x"30", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"66", x"22", x"00", x"66", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"78", x"7C", x"7E", x"7E", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"3F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7E", x"7C", x"7E", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"3F", x"3F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7F", x"7F", x"7F", x"7E", x"7E", x"7C", x"78", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"78", x"78", x"78", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1E", x"38", x"70", x"60", x"E0", x"C0", x"03", x"0F", x"1E", x"38", x"73", x"67", x"EE", x"CC", x"C1", x"C1", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"DC", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", 
															x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"E0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"3F", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"80", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FC", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"01", x"00", x"00", x"07", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"78", x"1C", x"0E", x"06", x"07", x"03", x"C0", x"F0", x"78", x"1C", x"CE", x"E6", x"77", x"33", x"83", x"83", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"3B", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", 
															x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C1", x"C1", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"DC", x"C0", x"E0", x"60", x"70", x"38", x"1E", x"0F", x"03", x"CC", x"EE", x"67", x"73", x"38", x"1E", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"3F", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"80", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FC", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"FF", x"FF", x"00", x"FF", x"FF", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"83", x"83", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", x"3B", x"03", x"07", x"06", x"0E", x"1C", x"78", x"F0", x"C0", x"33", x"77", x"E6", x"CE", x"1C", x"78", x"F0", x"C0", 
															x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", x"1B", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CB", x"F3", x"C3", x"C1", x"00", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"7F", x"55", x"55", x"5F", x"9B", x"00", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"C1", x"00", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"7F", x"00", x"00", x"00", x"9B", x"00", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"CF", x"EF", x"00", x"F0", x"FC", x"FE", x"00", x"EF", x"EF", x"EF", x"00", x"FE", x"FE", x"FE", x"00", x"00", x"7E", x"3E", x"1E", x"0E", x"06", x"02", x"00", x"FE", x"82", x"C6", x"EE", x"EE", x"C6", x"82", x"FE", x"EE", x"EE", x"00", x"11", x"11", x"00", x"EE", x"EE", x"00", x"00", x"EE", x"FF", x"FF", x"EE", x"EE", x"EE", x"00", x"FF", x"FF", x"C3", x"C3", x"C3", x"81", x"00", x"FF", x"81", x"C3", x"FF", x"FF", x"C3", x"81", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"F7", x"BB", x"FE", x"ED", x"DD", x"DD", x"FF", x"FF", x"08", x"44", x"01", x"13", x"B3", x"BB", x"BB", x"FB", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FC", x"0E", x"09", x"FF", x"01", x"FF", x"FE", x"FC", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"11", x"33", x"BB", x"BF", x"BF", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"08", x"44", x"01", x"13", x"B3", x"BB", x"BB", x"FF", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"99", x"B9", x"FD", x"FD", x"08", x"1D", x"12", x"20", x"01", x"00", x"00", x"00", x"07", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"A6", x"D0", x"98", x"04", x"00", x"00", x"00", x"F0", x"50", x"00", x"00", x"00", x"00", x"00", x"00", x"33", x"71", x"28", x"3F", x"71", x"40", x"80", x"01", x"0F", x"0F", x"17", x"00", x"00", x"00", x"00", x"00", x"E4", x"06", x"6D", x"68", x"96", x"8D", x"80", x"00", x"F8", x"F8", x"90", x"90", x"08", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"7E", x"00", x"00", x"00", x"00", x"00", x"3C", x"C2", x"86", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"02", x"7E", x"3E", x"1E", x"06", x"02", x"00", x"00", x"FE", x"86", x"CE", x"EE", x"E6", x"C2", x"82", x"FC", x"1E", x"0E", x"06", x"02", x"02", x"00", x"00", x"00", x"EE", x"EE", x"C6", x"C2", x"BE", x"C2", x"00", x"00", x"40", x"3E", x"1E", x"1E", x"0E", x"06", x"02", x"00", x"BE", x"C2", x"E6", x"EE", x"CE", x"86", x"C2", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"0E", x"00", x"00", x"00", x"00", x"3C", x"7E", x"1E", x"0E", x"00", x"00", x"00", x"3C", x"C2", x"86", x"EE", x"EE", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"B0", x"0E", x"7E", x"3E", x"0E", x"06", x"00", x"00", x"00", x"F2", x"86", x"CE", x"EE", x"E6", x"C2", x"8C", x"F0", x"06", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"C6", x"C2", x"BE", x"C2", x"00", x"00", x"00", x"00", x"30", x"3E", x"1E", x"0E", x"0E", x"06", x"02", x"00", x"CE", x"C2", x"E6", x"EE", x"8E", x"46", x"32", x"0E", x"00", x"00", x"00", x"00", x"02", x"06", x"0E", x"3E", x"00", x"00", x"00", x"02", x"06", x"0A", x"36", x"C6", x"00", x"00", x"3C", x"7E", x"1E", x"0E", x"06", x"02", x"00", x"3C", x"C2", x"86", x"EE", x"EE", x"C6", x"C2", x"00", x"00", x"00", x"00", x"40", x"20", x"30", x"1C", x"00", x"00", x"00", x"C0", x"A0", x"D0", x"CC", x"E2", x"7E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"8E", x"EE", x"E2", x"C4", x"C8", x"B0", x"C0", x"00", 
															x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BE", x"C2", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"0E", x"0E", x"06", x"02", x"02", x"00", x"00", x"E6", x"8E", x"CE", x"26", x"12", x"0E", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"E0", x"01", x"11", x"10", x"0E", x"EE", x"E0", x"00", x"0E", x"EF", x"FF", x"FE", x"EE", x"EE", x"E0", x"00", x"10", x"11", x"01", x"EE", x"EE", x"00", x"00", x"EE", x"FE", x"FF", x"EF", x"EE", x"EE", x"00", x"00", x"EE", x"0E", x"00", x"11", x"11", x"E0", x"EE", x"0E", x"00", x"E0", x"EE", x"FF", x"FF", x"EE", x"EE", x"0E", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"EE", x"00", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"EE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E1", x"E1", x"00", x"10", x"1E", x"0E", x"E0", x"E0", x"0F", x"0F", x"EE", x"FE", x"FE", x"EE", x"E0", x"E0", x"01", x"EF", x"EE", x"00", x"00", x"00", x"00", x"00", x"EF", x"EF", x"EE", x"00", x"00", x"00", x"00", x"00", x"0E", x"0E", x"00", x"11", x"F1", x"E0", x"0E", x"0E", x"E0", x"E0", x"EE", x"FF", x"FF", x"EE", x"0E", x"0E", x"00", x"00", x"00", x"00", x"0E", x"0E", x"E1", x"E1", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"00", x"EE", x"EE", x"00", x"10", x"10", x"01", x"EF", x"00", x"00", x"00", x"EE", x"FE", x"FE", x"EF", x"EF", 
															x"00", x"00", x"00", x"00", x"E0", x"E0", x"0E", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"00", x"10", x"1E", x"0E", x"E0", x"E0", x"00", x"00", x"EE", x"FE", x"FE", x"EE", x"E0", x"E0", x"00", x"00", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"F0", x"E1", x"0F", x"0E", x"00", x"00", x"EE", x"FE", x"FE", x"EF", x"0F", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"00", x"00", x"00", x"00", x"00", x"3C", x"C3", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"03", x"FF", x"FF", x"C3", x"C3", x"C1", x"80", x"00", x"FD", x"83", x"C3", x"FF", x"FF", x"C1", x"83", x"FC", 
															x"C3", x"C3", x"C3", x"C3", x"81", x"00", x"00", x"00", x"FF", x"FF", x"C3", x"C3", x"BD", x"C3", x"00", x"00", x"C0", x"FF", x"FF", x"C3", x"C3", x"83", x"01", x"00", x"BF", x"C1", x"C3", x"FF", x"FF", x"83", x"C1", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"0D", x"00", x"00", x"00", x"00", x"3C", x"FF", x"C3", x"C3", x"00", x"00", x"00", x"3C", x"C3", x"81", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"F0", x"0F", x"FF", x"F3", x"C3", x"C0", x"C0", x"80", x"00", x"F3", x"83", x"CF", x"FF", x"F1", x"C2", x"8C", x"F0", x"C3", x"C3", x"81", x"00", x"00", x"00", x"00", x"00", x"C3", x"C3", x"BD", x"C3", x"00", x"00", x"00", x"00", x"F0", x"FF", x"CF", x"83", x"03", x"03", x"01", x"00", x"CF", x"C1", x"F3", x"FF", x"8F", x"43", x"31", x"0F", 
															x"00", x"00", x"00", x"00", x"01", x"07", x"0F", x"3B", x"00", x"00", x"00", x"03", x"07", x"0B", x"33", x"C7", x"00", x"00", x"3C", x"FF", x"C3", x"C3", x"C3", x"C3", x"00", x"3C", x"C3", x"81", x"FF", x"FF", x"C3", x"C3", x"00", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"DC", x"00", x"00", x"00", x"C0", x"A0", x"D0", x"CC", x"E3", x"F3", x"C1", x"C0", x"C0", x"C0", x"80", x"00", x"00", x"8F", x"F9", x"F3", x"C4", x"C8", x"B0", x"C0", x"00", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BD", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"CF", x"83", x"03", x"03", x"03", x"01", x"00", x"00", x"F1", x"9F", x"CF", x"23", x"13", x"0D", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"00", x"00", x"00", x"00", x"00", x"3C", x"C3", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"03", x"FF", x"FC", x"00", x"03", x"FF", x"FC", x"00", x"FC", x"00", x"03", x"FC", x"03", x"FF", x"FF", x"FC", x"C3", x"00", x"3C", x"FF", x"C3", x"00", x"00", x"00", x"3C", x"C3", x"3C", x"FF", x"FF", x"C3", x"00", x"00", x"C0", x"FF", x"3F", x"00", x"C0", x"FF", x"3F", x"00", x"3F", x"00", x"C0", x"3F", x"C0", x"FF", x"FF", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"0C", x"00", x"00", x"00", x"00", x"3C", x"FF", x"C3", x"00", x"00", x"00", x"00", x"3C", x"C3", x"00", x"3C", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"00", x"00", x"00", x"00", x"00", x"80", x"40", x"30", x"0E", x"FC", x"F1", x"03", x"0E", x"FC", x"F0", x"00", x"F1", x"02", x"0D", x"F3", x"0F", x"FE", x"FC", x"F0", 
															x"3C", x"FF", x"C3", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"FF", x"C3", x"00", x"00", x"00", x"00", x"70", x"3F", x"8F", x"C0", x"70", x"3F", x"0F", x"00", x"8F", x"40", x"B0", x"CF", x"F0", x"7F", x"3F", x"0F", x"00", x"00", x"00", x"00", x"03", x"07", x"0C", x"38", x"00", x"00", x"00", x"03", x"04", x"08", x"33", x"C4", x"00", x"00", x"3C", x"FF", x"C3", x"00", x"3C", x"FF", x"00", x"3C", x"C3", x"00", x"3C", x"C3", x"3C", x"FF", x"00", x"00", x"00", x"00", x"C0", x"E0", x"30", x"1C", x"00", x"00", x"00", x"C0", x"20", x"10", x"CC", x"23", x"F3", x"C7", x"0C", x"38", x"F0", x"C0", x"00", x"00", x"0B", x"37", x"CF", x"3C", x"F8", x"F0", x"C0", x"00", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"CF", x"E3", x"30", x"1C", x"0F", x"03", x"00", x"00", x"D0", x"EC", x"F3", x"3C", x"1F", x"0F", x"03", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"F7", x"BB", x"FE", x"00", x"00", x"00", x"00", x"00", x"08", x"44", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"BB", x"FE", x"ED", x"DD", x"DD", x"FF", x"FF", x"00", x"44", x"01", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"ED", x"DD", x"DD", x"FF", x"FF", x"00", x"00", x"00", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"00", x"00", x"BB", x"FE", x"ED", x"DD", x"DD", x"FF", x"FF", x"00", x"44", x"01", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F7", x"BB", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"44", x"00", x"00", x"00", x"F7", x"BB", x"FE", x"ED", x"DD", x"00", x"00", x"00", x"08", x"44", x"01", x"13", x"33", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"F7", x"BB", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"44", x"FE", x"ED", x"DD", x"DD", x"FF", x"FF", x"00", x"00", x"01", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"00", x"DD", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"BB", x"BB", x"FB", x"00", x"00", x"00", x"00", x"00", x"FE", x"ED", x"DD", x"DD", x"FF", x"FF", x"00", x"00", x"01", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F7", x"BB", x"FE", x"00", x"00", x"00", x"00", x"00", x"08", x"44", x"01", x"00", x"F7", x"BB", x"FE", x"ED", x"DD", x"DD", x"FF", x"00", x"08", x"44", x"01", x"13", x"B3", x"BB", x"BB", x"00", x"00", x"00", x"00", x"00", x"F7", x"BB", x"FE", x"00", x"00", x"00", x"00", x"00", x"08", x"44", x"01", x"FD", x"DD", x"DD", x"FF", x"FF", x"00", x"00", x"00", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"00", x"00", 
															x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ED", x"DD", x"DD", x"FF", x"FF", x"00", x"00", x"00", x"13", x"B3", x"BB", x"BB", x"FB", x"00", x"00", x"00", x"00", x"7F", x"7F", x"00", x"F1", x"CB", x"CB", x"CB", x"7F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"00", x"95", x"55", x"55", x"55", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"00", x"F1", x"CB", x"CB", x"F3", x"7F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"00", x"95", x"55", x"55", x"5F", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"FB", x"CB", x"F3", x"7F", x"7F", x"7F", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"FE", x"D5", x"55", x"DF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF");
	
	constant SUPER_MARIO_CHR_ROM : CHR_ROM_ARRAY := (x"03", x"0F", x"1F", x"1F", x"1C", x"24", x"26", x"66", x"00", x"00", x"00", x"00", x"1F", x"3F", x"3F", x"7F", x"E0", x"C0", x"80", x"FC", x"80", x"C0", x"00", x"20", x"00", x"20", x"60", x"00", x"F0", x"FC", x"FE", x"FE", x"60", x"70", x"18", x"07", x"0F", x"1F", x"3F", x"7F", x"7F", x"7F", x"1F", x"07", x"00", x"1E", x"3F", x"7F", x"FC", x"7C", x"00", x"00", x"E0", x"F0", x"F8", x"F8", x"FC", x"FC", x"F8", x"C0", x"C2", x"67", x"2F", x"37", x"7F", x"7F", x"FF", x"FF", x"07", x"07", x"0F", x"0F", x"7F", x"7E", x"FC", x"F0", x"F8", x"F8", x"F0", x"70", x"FD", x"FE", x"B4", x"F8", x"F8", x"F9", x"FB", x"FF", x"37", x"36", x"5C", x"00", x"00", x"01", x"03", x"1F", x"1F", x"3F", x"FF", x"FF", x"FC", x"70", x"70", x"38", x"08", x"24", x"E3", x"F0", x"F8", x"70", x"70", x"38", x"FF", x"FF", x"FF", x"1F", x"00", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"01", x"07", x"0F", x"0F", x"0E", x"12", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"00", x"00", x"F0", x"E0", x"C0", x"FE", x"40", x"60", x"00", x"00", x"00", x"10", x"30", x"00", x"F8", x"FE", x"13", x"33", x"30", x"18", x"04", x"0F", x"1F", x"1F", x"1F", x"3F", x"3F", x"1F", x"07", x"08", x"17", x"17", x"00", x"10", x"7E", x"3E", x"00", x"00", x"C0", x"E0", x"FF", x"FF", x"FE", x"FE", x"FC", x"E0", x"40", x"A0", x"3F", x"3F", x"3F", x"1F", x"1F", x"1F", x"1F", x"1F", x"37", x"27", x"23", x"03", x"01", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F8", x"F8", x"F8", x"F8", x"F8", x"CC", x"FF", x"FF", x"FF", x"FF", x"70", x"00", x"08", x"FF", x"FF", x"FF", x"FE", x"F0", x"C0", x"80", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"C0", x"80", x"00", x"FC", x"FC", x"F8", x"78", x"78", x"78", x"7E", x"7E", x"10", x"60", x"80", x"00", x"78", x"78", x"7E", x"7E", 
															x"00", x"03", x"0F", x"1F", x"1F", x"1C", x"24", x"26", x"00", x"00", x"00", x"00", x"00", x"1F", x"3F", x"3F", x"00", x"E0", x"C0", x"80", x"FC", x"80", x"C0", x"00", x"00", x"00", x"20", x"60", x"00", x"F0", x"FC", x"FE", x"66", x"60", x"30", x"18", x"0F", x"1F", x"3F", x"3F", x"7F", x"7F", x"3F", x"1F", x"00", x"16", x"2F", x"2F", x"20", x"FC", x"7C", x"00", x"00", x"E0", x"E0", x"F0", x"FE", x"FC", x"FC", x"F8", x"C0", x"60", x"20", x"30", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"1F", x"2F", x"2F", x"2F", x"0F", x"07", x"03", x"00", x"00", x"F0", x"90", x"00", x"08", x"0C", x"1C", x"FC", x"F8", x"10", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"E0", x"0F", x"0F", x"07", x"07", x"07", x"0F", x"0F", x"03", x"01", x"03", x"01", x"04", x"07", x"0F", x"0F", x"03", x"F8", x"F0", x"E0", x"F0", x"B0", x"80", x"E0", x"E0", x"F8", x"F0", x"E0", x"70", x"B0", x"80", x"E0", x"E0", 
															x"03", x"3F", x"7F", x"19", x"09", x"09", x"28", x"5C", x"00", x"30", x"70", x"7F", x"FF", x"FF", x"F7", x"F3", x"F8", x"E0", x"E0", x"FC", x"26", x"30", x"80", x"10", x"00", x"18", x"10", x"00", x"F8", x"F8", x"FE", x"FF", x"3E", x"1E", x"3F", x"38", x"30", x"30", x"00", x"3A", x"E7", x"0F", x"0F", x"1F", x"1F", x"1F", x"0F", x"07", x"78", x"1E", x"80", x"FE", x"7E", x"7E", x"7F", x"7F", x"FF", x"FE", x"FC", x"C6", x"8E", x"EE", x"FF", x"FF", x"3C", x"3F", x"1F", x"0F", x"07", x"3F", x"21", x"20", x"03", x"00", x"00", x"0E", x"07", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FC", x"70", x"FF", x"7F", x"3F", x"0E", x"C0", x"C0", x"E0", x"E0", x"0F", x"9F", x"CF", x"FF", x"7F", x"3F", x"1E", x"0E", x"00", x"80", x"C8", x"FE", x"7F", x"3F", x"1E", x"0E", x"20", x"C0", x"80", x"80", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"03", x"0F", x"1F", x"1F", x"1C", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"3F", x"00", x"04", x"E6", x"E0", x"FF", x"FF", x"8F", x"83", x"0E", x"1F", x"1F", x"1F", x"1F", x"03", x"FF", x"FF", x"26", x"26", x"60", x"78", x"18", x"0F", x"7F", x"FF", x"3F", x"3F", x"7F", x"7F", x"1F", x"00", x"7E", x"FF", x"01", x"21", x"FE", x"7A", x"06", x"FE", x"FC", x"FC", x"FF", x"FF", x"FE", x"FE", x"FE", x"DE", x"5C", x"6C", x"FF", x"CF", x"87", x"07", x"07", x"0F", x"1F", x"1F", x"FF", x"FF", x"FE", x"FC", x"F8", x"B0", x"60", x"00", x"F8", x"F8", x"F0", x"B8", x"F8", x"F9", x"FB", x"FF", x"28", x"30", x"18", x"40", x"00", x"01", x"03", x"0F", x"1F", x"FF", x"FF", x"FF", x"FF", x"FE", x"C0", x"80", x"10", x"EC", x"E3", x"E0", x"E0", x"E0", x"C0", x"80", x"FF", x"FF", x"FF", x"3F", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", 
															x"13", x"33", x"30", x"18", x"04", x"0F", x"1F", x"1F", x"1F", x"3F", x"3F", x"1F", x"07", x"09", x"13", x"17", x"00", x"10", x"7E", x"30", x"E0", x"F0", x"F0", x"E0", x"FF", x"FF", x"FE", x"FF", x"FE", x"FC", x"F8", x"E0", x"1F", x"1F", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"17", x"17", x"03", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F8", x"F8", x"B8", x"F8", x"F8", x"F8", x"D0", x"90", x"18", x"08", x"40", x"00", x"00", x"00", x"3F", x"FF", x"FF", x"FF", x"F6", x"C6", x"84", x"00", x"30", x"F0", x"F0", x"F1", x"F6", x"C6", x"84", x"00", x"F0", x"E0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"3F", x"3F", x"1F", x"0F", x"0F", x"1F", x"1F", x"1F", x"3F", x"3E", x"7C", x"78", x"F0", x"E0", x"F0", x"F0", x"F8", x"F8", x"B8", x"F8", x"F8", x"F0", x"B0", x"90", x"18", x"08", x"40", x"00", x"00", x"00", 
															x"E0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F8", x"F0", x"C0", x"E0", x"FC", x"FE", x"FF", x"7F", x"03", x"00", x"1F", x"1F", x"1F", x"3F", x"3E", x"3C", x"38", x"18", x"00", x"00", x"10", x"38", x"3E", x"3C", x"38", x"18", x"00", x"03", x"07", x"07", x"0A", x"0B", x"0C", x"00", x"00", x"00", x"00", x"07", x"0F", x"0F", x"0F", x"03", x"00", x"E0", x"FC", x"20", x"20", x"10", x"3C", x"00", x"00", x"00", x"00", x"F0", x"FC", x"FE", x"FC", x"F8", x"07", x"07", x"07", x"1F", x"1F", x"3E", x"21", x"01", x"07", x"0F", x"1B", x"18", x"10", x"30", x"21", x"01", x"E0", x"E0", x"E0", x"F0", x"F0", x"E0", x"C0", x"E0", x"A8", x"FC", x"F8", x"00", x"00", x"00", x"C0", x"E0", x"07", x"0F", x"0E", x"14", x"16", x"18", x"00", x"3F", x"00", x"00", x"0F", x"1F", x"1F", x"1F", x"07", x"3C", x"C0", x"F8", x"40", x"40", x"20", x"78", x"00", x"C0", x"00", x"00", x"E0", x"F8", x"FC", x"F8", x"F0", x"C0", 
															x"3F", x"0E", x"0F", x"1F", x"3F", x"7C", x"70", x"38", x"FC", x"ED", x"C0", x"00", x"00", x"60", x"70", x"38", x"F0", x"F8", x"E4", x"FC", x"FC", x"7C", x"00", x"00", x"7E", x"1E", x"04", x"0C", x"0C", x"0C", x"00", x"00", x"07", x"0F", x"0E", x"14", x"16", x"18", x"00", x"0F", x"00", x"00", x"0F", x"1F", x"1F", x"1F", x"07", x"0D", x"1F", x"1F", x"1F", x"1C", x"0C", x"07", x"07", x"07", x"1E", x"1C", x"1E", x"0F", x"07", x"00", x"07", x"07", x"E0", x"60", x"F0", x"70", x"E0", x"E0", x"F0", x"80", x"60", x"90", x"00", x"80", x"00", x"E0", x"F0", x"80", x"07", x"1F", x"3F", x"12", x"13", x"08", x"1F", x"31", x"00", x"10", x"3F", x"7F", x"7F", x"3F", x"03", x"0F", x"C0", x"F0", x"40", x"00", x"30", x"18", x"C0", x"F8", x"00", x"00", x"E0", x"F8", x"FC", x"F8", x"B0", x"38", x"31", x"39", x"1F", x"1F", x"0F", x"5F", x"7E", x"3C", x"1F", x"07", x"00", x"0E", x"0F", x"53", x"7C", x"3C", 
															x"F8", x"F8", x"F0", x"E0", x"E0", x"C0", x"00", x"00", x"F8", x"F8", x"F0", x"00", x"00", x"80", x"00", x"00", x"00", x"E0", x"FC", x"27", x"27", x"11", x"3E", x"04", x"07", x"07", x"03", x"F7", x"FF", x"FF", x"FE", x"FC", x"3F", x"7F", x"3F", x"0F", x"1F", x"3F", x"7F", x"4F", x"3E", x"7F", x"FF", x"E2", x"50", x"38", x"70", x"40", x"F8", x"F9", x"F9", x"B7", x"FF", x"FF", x"E0", x"00", x"E8", x"71", x"01", x"4B", x"03", x"03", x"00", x"00", x"07", x"07", x"0F", x"3F", x"3F", x"3F", x"26", x"04", x"05", x"03", x"01", x"30", x"30", x"30", x"26", x"04", x"F0", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"FE", x"FC", x"E0", x"00", x"00", x"00", x"00", x"00", x"07", x"07", x"0F", x"1F", x"3F", x"0F", x"1C", x"18", x"05", x"03", x"01", x"10", x"30", x"0C", x"1C", x"18", x"E0", x"E0", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"C0", x"E0", x"F0", x"78", x"18", x"08", x"00", x"00", 
															x"07", x"0F", x"1F", x"0F", x"3F", x"0F", x"1C", x"18", x"07", x"0F", x"3E", x"7C", x"30", x"0C", x"1C", x"18", x"E0", x"E0", x"E0", x"40", x"C0", x"80", x"00", x"00", x"60", x"60", x"60", x"80", x"00", x"00", x"00", x"00", x"7F", x"FF", x"FF", x"FB", x"0F", x"0F", x"0F", x"1F", x"73", x"F3", x"F0", x"F4", x"F0", x"F0", x"70", x"60", x"3F", x"7E", x"7C", x"7C", x"3C", x"3C", x"FC", x"FC", x"00", x"00", x"00", x"00", x"3C", x"3C", x"FC", x"FC", x"60", x"70", x"18", x"08", x"0F", x"1F", x"3F", x"7F", x"7F", x"7F", x"1F", x"07", x"0B", x"1B", x"3B", x"7B", x"FC", x"7C", x"00", x"20", x"F0", x"F8", x"FC", x"FE", x"FC", x"FC", x"F8", x"E0", x"D0", x"D8", x"DC", x"DE", x"0B", x"0F", x"1F", x"1E", x"3C", x"3C", x"3C", x"7C", x"C4", x"E0", x"E0", x"40", x"00", x"3C", x"3C", x"7C", x"1F", x"3F", x"0D", x"07", x"0F", x"0E", x"1C", x"3C", x"1D", x"3C", x"3A", x"38", x"30", x"00", x"1C", x"3C", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"22", x"55", x"55", x"55", x"55", x"55", x"77", x"22", x"00", x"07", x"1F", x"FF", x"07", x"1F", x"0F", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"76", x"00", x"00", x"CF", x"07", x"7F", x"00", x"00", x"00", x"20", x"F8", x"FF", x"C3", x"FD", x"FE", x"F0", x"40", x"00", x"00", x"3C", x"FC", x"FE", x"E0", x"00", x"00", x"40", x"E0", x"40", x"40", x"41", x"41", x"4F", x"47", x"40", x"E0", x"40", x"3F", x"3E", x"3E", x"30", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"C0", x"00", x"00", x"00", x"F8", x"F8", x"F8", x"18", x"38", x"43", x"46", x"44", x"40", x"40", x"40", x"40", x"40", x"3C", x"39", x"3B", x"3F", x"00", x"00", x"00", x"00", x"80", x"C0", x"40", x"00", x"00", x"00", x"00", x"00", x"78", x"38", x"B8", x"F8", x"00", x"00", x"00", x"00", 
															x"31", x"30", x"38", x"7C", x"7F", x"FF", x"FF", x"FB", x"3F", x"3F", x"0F", x"77", x"77", x"F7", x"F7", x"F7", x"10", x"7E", x"3E", x"00", x"1E", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FA", x"FA", x"F3", x"E7", x"FF", x"FF", x"E3", x"C3", x"87", x"48", x"3C", x"FC", x"F0", x"F8", x"FC", x"7C", x"78", x"38", x"3C", x"FC", x"00", x"FF", x"C3", x"83", x"83", x"FF", x"FF", x"FF", x"FF", x"00", x"C3", x"81", x"81", x"C3", x"FF", x"00", x"1F", x"1F", x"0F", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"FB", x"FF", x"FF", x"FE", x"3E", x"0C", x"04", x"00", x"0B", x"1F", x"1F", x"1E", x"3E", x"0C", x"04", x"1F", x"1F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FB", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"03", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", 
															x"00", x"18", x"3C", x"7E", x"6E", x"DF", x"DF", x"DF", x"00", x"18", x"3C", x"7E", x"76", x"FB", x"FB", x"FB", x"00", x"18", x"18", x"3C", x"3C", x"3C", x"3C", x"1C", x"00", x"10", x"10", x"20", x"20", x"20", x"20", x"20", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"08", x"08", x"04", x"04", x"04", x"04", x"04", x"00", x"10", x"10", x"38", x"38", x"38", x"38", x"38", x"3C", x"7E", x"77", x"FB", x"9F", x"5F", x"8E", x"20", x"00", x"18", x"3C", x"0E", x"0E", x"04", x"00", x"00", x"5C", x"2E", x"8F", x"3F", x"7B", x"77", x"7E", x"3C", x"00", x"00", x"04", x"06", x"1E", x"3C", x"18", x"00", x"13", x"4F", x"3F", x"BF", x"3F", x"7A", x"F8", x"F8", x"00", x"00", x"01", x"0A", x"17", x"0F", x"2F", x"1F", x"00", x"08", x"05", x"0F", x"2F", x"1D", x"1C", x"3C", x"00", x"00", x"00", x"00", x"05", x"07", x"0F", x"07", 
															x"00", x"00", x"00", x"00", x"02", x"0B", x"07", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"08", x"04", x"04", x"00", x"60", x"F0", x"F8", x"7C", x"3E", x"7E", x"7F", x"02", x"02", x"02", x"05", x"71", x"7F", x"7F", x"7F", x"3F", x"5F", x"7F", x"3E", x"0E", x"0A", x"51", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"1F", x"02", x"02", x"00", x"01", x"13", x"3F", x"7F", x"7F", x"3F", x"7F", x"7F", x"FE", x"EC", x"CA", x"51", x"20", x"00", x"40", x"60", x"70", x"73", x"27", x"0F", x"1F", x"00", x"40", x"63", x"77", x"7C", x"38", x"F8", x"E4", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"1F", x"00", x"00", x"03", x"07", x"0C", x"18", x"F8", x"E4", x"7F", x"7F", x"3F", x"3F", x"1F", x"1F", x"0F", x"07", x"03", x"44", x"28", x"10", x"08", x"04", x"03", x"04", 
															x"03", x"07", x"0F", x"1F", x"3F", x"77", x"77", x"F5", x"03", x"07", x"0F", x"1F", x"27", x"7B", x"78", x"FB", x"C0", x"E0", x"F0", x"F8", x"FC", x"EE", x"EE", x"AF", x"C0", x"E0", x"F0", x"F8", x"E4", x"DE", x"1E", x"DF", x"F1", x"FF", x"78", x"00", x"00", x"18", x"1C", x"0E", x"FF", x"FF", x"7F", x"0F", x"0F", x"07", x"03", x"00", x"8F", x"FF", x"1E", x"00", x"0C", x"3E", x"7E", x"7C", x"FF", x"FF", x"FE", x"F0", x"F0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"24", x"24", x"18", x"00", x"00", x"00", x"02", x"41", x"41", x"61", x"33", x"06", x"3C", x"3C", x"7E", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"7F", x"FF", x"03", x"07", x"0F", x"1F", x"3F", x"63", x"41", x"C1", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FE", x"FF", x"C0", x"80", x"00", x"00", x"8C", x"FE", x"FE", x"F3", 
															x"FF", x"FF", x"FF", x"78", x"00", x"00", x"00", x"00", x"C1", x"E3", x"FF", x"47", x"0F", x"0F", x"0F", x"07", x"FF", x"FF", x"FF", x"1E", x"00", x"20", x"20", x"40", x"F1", x"F9", x"FF", x"E2", x"F0", x"F0", x"F0", x"E0", x"16", x"1F", x"3F", x"7F", x"3D", x"1D", x"3F", x"1F", x"16", x"1F", x"00", x"00", x"05", x"0D", x"3F", x"1F", x"80", x"80", x"C0", x"E0", x"F0", x"F0", x"F0", x"F8", x"80", x"80", x"00", x"00", x"00", x"A0", x"A0", x"E0", x"3C", x"FA", x"B1", x"72", x"F2", x"DB", x"DF", x"5F", x"00", x"04", x"4E", x"8C", x"0C", x"7F", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"06", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", x"00", x"7C", x"D6", x"92", x"BA", x"EE", x"FE", x"38", x"FF", x"83", x"29", x"6D", x"45", x"11", x"01", x"C7", 
															x"00", x"15", x"3F", x"62", x"5F", x"FF", x"9F", x"7D", x"08", x"08", x"02", x"1F", x"22", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"2F", x"1E", x"2F", x"2F", x"2F", x"15", x"0D", x"0E", x"10", x"1E", x"10", x"50", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"1C", x"3E", x"7F", x"FF", x"FF", x"FE", x"7C", x"38", x"1C", x"2A", x"77", x"EE", x"DD", x"AA", x"74", x"28", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"00", x"EF", x"EF", x"EF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"00", x"EF", x"EF", x"EF", x"00", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7F", x"5F", x"7F", x"7F", x"7F", x"7F", x"7F", 
															x"68", x"4E", x"E0", x"E0", x"E0", x"F0", x"F8", x"FC", x"B8", x"9E", x"80", x"C0", x"E0", x"F0", x"F8", x"7C", x"3F", x"5C", x"39", x"3B", x"BB", x"F9", x"FC", x"FE", x"00", x"23", x"57", x"4F", x"57", x"27", x"C3", x"21", x"C0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"30", x"70", x"70", x"F0", x"E0", x"C0", x"00", x"FE", x"FC", x"61", x"0F", x"FF", x"FE", x"F0", x"E0", x"13", x"0F", x"1E", x"F0", x"FC", x"F8", x"F0", x"E0", x"6E", x"40", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"BE", x"90", x"80", x"C0", x"C0", x"80", x"00", x"00", x"01", x"01", x"03", x"03", x"07", x"7F", x"7F", x"3F", x"01", x"01", x"03", x"03", x"07", x"7F", x"7D", x"3D", x"06", x"07", x"3F", x"3C", x"19", x"7B", x"7F", x"3F", x"06", x"04", x"30", x"23", x"06", x"64", x"60", x"00", x"3F", x"7F", x"7F", x"1F", x"3F", x"3F", x"07", x"06", x"00", x"60", x"60", x"00", x"20", x"30", x"04", x"06", 
															x"03", x"07", x"0F", x"0F", x"0F", x"0F", x"07", x"03", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"F8", x"F8", x"F8", x"A0", x"E1", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"40", x"01", x"03", x"03", x"03", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"0F", x"07", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"F8", x"F8", x"FF", x"FE", x"F0", x"C0", x"E0", x"FE", x"FF", x"7F", x"03", x"02", x"00", x"00", x"01", x"0F", x"0F", x"1F", x"39", x"33", x"37", x"7F", x"01", x"0D", x"08", x"00", x"36", x"2C", x"08", x"60", x"7F", x"3F", x"3F", x"3F", x"1F", x"0F", x"0F", x"01", x"60", x"00", x"20", x"30", x"00", x"08", x"0D", x"01", x"00", x"00", x"03", x"03", x"47", x"67", x"77", x"77", x"01", x"01", x"03", x"43", x"67", x"77", x"7B", x"78", x"00", x"00", x"00", x"00", x"88", x"98", x"F8", x"F0", x"00", x"00", x"80", x"84", x"CC", x"DC", x"BC", x"3C", 
															x"7E", x"7F", x"FF", x"1F", x"07", x"30", x"1C", x"0C", x"33", x"07", x"07", x"E3", x"38", x"3F", x"1C", x"0C", x"7E", x"38", x"F6", x"ED", x"DF", x"38", x"70", x"60", x"98", x"C7", x"C8", x"92", x"30", x"F8", x"70", x"60", x"00", x"00", x"00", x"03", x"03", x"47", x"67", x"77", x"00", x"01", x"01", x"03", x"43", x"67", x"77", x"7B", x"00", x"00", x"00", x"00", x"00", x"88", x"98", x"F8", x"00", x"00", x"00", x"80", x"84", x"CC", x"DC", x"BC", x"77", x"7E", x"7F", x"FF", x"1F", x"07", x"70", x"F0", x"78", x"33", x"07", x"07", x"E3", x"38", x"7F", x"F0", x"F0", x"7E", x"38", x"F6", x"ED", x"DF", x"38", x"3C", x"3C", x"98", x"C7", x"C8", x"92", x"30", x"F8", x"3C", x"03", x"07", x"0A", x"1A", x"1C", x"1E", x"0B", x"08", x"00", x"10", x"7F", x"7F", x"7F", x"1F", x"0F", x"0F", x"1C", x"3F", x"3F", x"3D", x"3F", x"1F", x"00", x"00", x"03", x"33", x"39", x"3A", x"38", x"18", x"00", x"00", 
															x"00", x"00", x"04", x"4C", x"4E", x"4E", x"46", x"6F", x"10", x"38", x"3C", x"74", x"76", x"76", x"7E", x"7D", x"00", x"1F", x"3F", x"3F", x"4F", x"5F", x"7F", x"7F", x"00", x"00", x"11", x"0A", x"34", x"2A", x"51", x"20", x"7F", x"67", x"A3", x"B0", x"D8", x"DE", x"DC", x"C8", x"7F", x"67", x"63", x"70", x"38", x"3E", x"7C", x"B8", x"7F", x"7F", x"7F", x"1F", x"47", x"70", x"70", x"39", x"51", x"0A", x"04", x"EA", x"79", x"7F", x"70", x"39", x"E8", x"E8", x"E0", x"C0", x"10", x"70", x"E0", x"C0", x"58", x"38", x"10", x"30", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"20", x"66", x"66", x"66", x"62", x"00", x"08", x"1C", x"3C", x"7A", x"7A", x"7A", x"7E", x"00", x"00", x"1F", x"3F", x"7F", x"4F", x"5F", x"7F", x"00", x"00", x"00", x"11", x"0A", x"34", x"2A", x"51", x"77", x"7F", x"3F", x"B7", x"B3", x"DB", x"DA", x"D8", x"7F", x"7D", x"3F", x"37", x"33", x"3B", x"3A", x"78", 
															x"7F", x"7F", x"7F", x"7F", x"1F", x"07", x"70", x"F0", x"20", x"51", x"0A", x"04", x"EA", x"39", x"7F", x"F0", x"CC", x"E8", x"E8", x"E0", x"C0", x"18", x"7C", x"3E", x"BC", x"58", x"38", x"10", x"30", x"F8", x"FC", x"3E", x"03", x"0F", x"1F", x"3F", x"3B", x"3F", x"7F", x"7F", x"00", x"00", x"00", x"06", x"0E", x"0C", x"00", x"00", x"80", x"F0", x"F8", x"FC", x"FE", x"FE", x"FF", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"18", x"7F", x"7F", x"7F", x"7F", x"FF", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"F8", x"3E", x"3B", x"18", x"FE", x"FB", x"FF", x"FF", x"F6", x"E0", x"C0", x"00", x"10", x"14", x"10", x"10", x"38", x"78", x"F8", x"30", x"00", x"03", x"0F", x"1F", x"3F", x"3B", x"3F", x"7F", x"00", x"00", x"00", x"00", x"06", x"0E", x"0C", x"00", x"00", x"C0", x"F0", x"F8", x"FC", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", 
															x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"F8", x"7E", x"F3", x"FE", x"FE", x"FB", x"FF", x"FF", x"F6", x"E0", x"C0", x"18", x"10", x"14", x"10", x"10", x"38", x"7C", x"DE", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"08", x"00", x"0D", x"1E", x"1E", x"1E", x"1F", x"0F", x"07", x"78", x"F0", x"F8", x"E4", x"C0", x"CA", x"CA", x"C0", x"78", x"F0", x"00", x"1A", x"3F", x"35", x"35", x"3F", x"0F", x"1F", x"9F", x"FF", x"FF", x"7F", x"74", x"20", x"00", x"00", x"80", x"E0", x"E0", x"70", x"73", x"21", x"E4", x"FF", x"FE", x"FC", x"9C", x"1E", x"00", x"00", x"1A", x"07", x"0C", x"18", x"78", x"FE", x"FC", x"F0", x"00", x"01", x"03", x"03", x"07", x"03", x"01", x"00", x"00", x"01", x"02", x"00", x"38", x"7C", x"7E", x"3F", x"00", x"5F", x"7F", x"7F", x"3F", x"3F", x"14", x"00", x"3F", x"40", x"60", x"60", x"20", x"30", x"13", x"01", 
															x"C0", x"E0", x"F0", x"30", x"38", x"3C", x"3C", x"FC", x"C0", x"E0", x"30", x"D0", x"D0", x"D0", x"D0", x"00", x"07", x"0F", x"1F", x"22", x"20", x"25", x"25", x"1F", x"07", x"0F", x"02", x"1D", x"1F", x"1A", x"1A", x"02", x"FE", x"FE", x"7E", x"3A", x"02", x"01", x"41", x"41", x"38", x"7C", x"FC", x"FC", x"FC", x"FE", x"BE", x"BE", x"1F", x"3F", x"7E", x"5C", x"40", x"80", x"82", x"82", x"1C", x"3E", x"3F", x"3F", x"3F", x"7F", x"7D", x"7D", x"82", x"80", x"A0", x"44", x"43", x"40", x"21", x"1E", x"7D", x"7F", x"5F", x"3B", x"3C", x"3F", x"1E", x"00", x"1C", x"3F", x"3E", x"3C", x"40", x"80", x"82", x"82", x"1C", x"3E", x"3F", x"1F", x"3F", x"7F", x"7D", x"7D", x"00", x"00", x"80", x"80", x"92", x"9D", x"C7", x"EF", x"00", x"00", x"00", x"60", x"62", x"65", x"3F", x"1F", x"00", x"23", x"33", x"3F", x"3F", x"7F", x"7F", x"7F", x"70", x"3C", x"3C", x"18", x"00", x"00", x"02", x"07", 
															x"FE", x"F8", x"A0", x"00", x"00", x"00", x"80", x"80", x"CF", x"7A", x"5A", x"10", x"00", x"00", x"C0", x"80", x"7E", x"7F", x"7D", x"3F", x"1E", x"8F", x"8F", x"19", x"85", x"84", x"86", x"C6", x"E7", x"73", x"73", x"E1", x"E0", x"0E", x"73", x"F3", x"F9", x"F9", x"F8", x"70", x"80", x"4E", x"77", x"F3", x"FB", x"F9", x"FA", x"78", x"0E", x"66", x"E2", x"F6", x"FF", x"FF", x"1F", x"98", x"11", x"39", x"7D", x"39", x"00", x"00", x"E0", x"E7", x"00", x"00", x"00", x"04", x"0F", x"0F", x"1F", x"07", x"00", x"00", x"07", x"07", x"16", x"10", x"00", x"38", x"F3", x"E7", x"EE", x"EC", x"CD", x"CF", x"CF", x"DF", x"CF", x"1F", x"17", x"10", x"33", x"30", x"30", x"20", x"27", x"3F", x"3F", x"78", x"3C", x"1F", x"1F", x"73", x"38", x"30", x"40", x"C7", x"07", x"66", x"E0", x"6C", x"9F", x"3E", x"7C", x"FC", x"F8", x"F8", x"C0", x"40", x"60", x"C0", x"80", x"04", x"9E", x"FF", x"F0", x"F8", 
															x"7F", x"7E", x"78", x"01", x"07", x"1F", x"3C", x"7C", x"24", x"01", x"07", x"FE", x"FF", x"7F", x"3F", x"7F", x"FC", x"F8", x"A0", x"FE", x"FC", x"F0", x"80", x"00", x"CF", x"7A", x"0A", x"FE", x"FC", x"00", x"00", x"00", x"7E", x"7F", x"7F", x"3F", x"1F", x"8F", x"8F", x"18", x"85", x"86", x"83", x"C3", x"E1", x"70", x"70", x"E0", x"9F", x"3E", x"7C", x"F8", x"F8", x"3C", x"18", x"F8", x"60", x"C0", x"80", x"00", x"98", x"FC", x"FE", x"FF", x"7F", x"7F", x"78", x"01", x"07", x"13", x"F1", x"03", x"24", x"00", x"07", x"FE", x"FF", x"7F", x"FF", x"03", x"00", x"00", x"1C", x"1D", x"1B", x"C3", x"E3", x"E1", x"03", x"0F", x"23", x"62", x"64", x"3C", x"1C", x"1E", x"E0", x"CD", x"1D", x"4F", x"EE", x"FF", x"3F", x"3F", x"1F", x"3D", x"6D", x"4F", x"EE", x"F3", x"20", x"03", x"3F", x"3F", x"00", x"00", x"70", x"B8", x"FC", x"FC", x"07", x"07", x"1F", x"3F", x"0F", x"47", x"03", x"00", 
															x"07", x"0F", x"1F", x"3F", x"3E", x"7C", x"78", x"78", x"00", x"00", x"03", x"07", x"0F", x"0F", x"1F", x"1F", x"3F", x"5C", x"39", x"3B", x"BF", x"FF", x"FE", x"FE", x"00", x"23", x"57", x"4F", x"57", x"2F", x"DF", x"21", x"C0", x"C0", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"FE", x"FC", x"61", x"0F", x"7F", x"3F", x"1F", x"1E", x"23", x"0F", x"1E", x"F0", x"1C", x"3F", x"1F", x"1E", x"F0", x"78", x"E4", x"C8", x"CC", x"BE", x"BE", x"3E", x"00", x"80", x"18", x"30", x"34", x"FE", x"FE", x"FE", x"00", x"01", x"00", x"07", x"07", x"07", x"07", x"1F", x"00", x"00", x"01", x"04", x"06", x"06", x"07", x"07", x"00", x"00", x"0F", x"3F", x"3F", x"0F", x"00", x"00", x"0F", x"3F", x"7F", x"F8", x"F8", x"7F", x"3F", x"0F", x"78", x"7C", x"7E", x"7F", x"3F", x"3F", x"1B", x"09", x"1F", x"1F", x"1F", x"0B", x"01", x"01", x"00", x"00", 
															x"0C", x"00", x"00", x"00", x"07", x"7F", x"7C", x"00", x"03", x"1F", x"3F", x"3F", x"78", x"00", x"03", x"FF", x"01", x"E1", x"71", x"79", x"3D", x"3D", x"1F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"1F", x"1B", x"36", x"30", x"7F", x"3F", x"23", x"27", x"1F", x"07", x"0F", x"1F", x"7F", x"3F", x"F8", x"F8", x"F8", x"B8", x"18", x"D8", x"D8", x"B8", x"E0", x"80", x"80", x"40", x"E0", x"E0", x"E0", x"C0", x"01", x"02", x"04", x"04", x"08", x"08", x"10", x"10", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"1F", x"00", x"0F", x"13", x"0D", x"0D", x"13", x"0C", x"20", x"1F", x"10", x"0C", x"12", x"12", x"2C", x"3F", x"3F", x"00", x"24", x"00", x"24", x"00", x"04", x"00", x"00", x"37", x"36", x"36", x"36", x"16", x"16", x"12", x"02", x"0F", x"41", x"00", x"88", x"00", x"44", x"00", x"00", x"10", x"7E", x"FF", x"FF", x"F6", x"76", x"3A", x"1A", 
															x"38", x"7C", x"FE", x"FE", x"3B", x"03", x"03", x"03", x"00", x"00", x"38", x"04", x"00", x"00", x"00", x"00", x"03", x"33", x"7B", x"7F", x"FF", x"FB", x"03", x"03", x"00", x"00", x"00", x"38", x"40", x"00", x"00", x"00", x"DC", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"FC", x"A0", x"80", x"80", x"00", x"00", x"00", x"00", x"3F", x"5F", x"3F", x"3F", x"BB", x"F8", x"FE", x"FE", x"07", x"27", x"57", x"4F", x"57", x"27", x"C1", x"21", x"1F", x"0F", x"0F", x"1F", x"1F", x"1E", x"38", x"30", x"1D", x"0F", x"0F", x"1F", x"1F", x"1E", x"38", x"30", x"00", x"20", x"60", x"60", x"70", x"F0", x"F8", x"F8", x"00", x"00", x"38", x"10", x"4C", x"18", x"86", x"24", x"F8", x"FC", x"FC", x"7E", x"7E", x"3E", x"1F", x"07", x"00", x"42", x"0A", x"40", x"10", x"02", x"08", x"02", x"00", x"C0", x"70", x"B8", x"F4", x"F2", x"F5", x"7B", x"00", x"00", x"80", x"40", x"08", x"0C", x"0A", x"84", 
															x"00", x"DF", x"10", x"FF", x"DF", x"FF", x"FF", x"F9", x"00", x"00", x"CF", x"20", x"20", x"20", x"26", x"2E", x"1F", x"1F", x"3E", x"FC", x"F8", x"F0", x"C0", x"00", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"F8", x"FC", x"FE", x"FF", x"FF", x"DF", x"DF", x"00", x"2F", x"23", x"21", x"20", x"20", x"00", x"00", x"00", x"C1", x"F1", x"79", x"7D", x"3D", x"3F", x"1F", x"03", x"C1", x"B1", x"59", x"6D", x"35", x"3B", x"1F", x"03", x"02", x"06", x"0E", x"0E", x"1E", x"1E", x"3E", x"3E", x"00", x"02", x"00", x"08", x"02", x"00", x"28", x"00", x"3E", x"3E", x"3E", x"3E", x"1E", x"1E", x"0E", x"02", x"04", x"10", x"02", x"10", x"04", x"00", x"0A", x"00", x"C1", x"F1", x"79", x"7D", x"3D", x"3F", x"1F", x"03", x"C1", x"B1", x"59", x"6D", x"35", x"3B", x"1F", x"03", x"7C", x"00", x"00", x"FF", x"C3", x"7F", x"1F", x"03", x"00", x"0F", x"1F", x"FF", x"FC", x"63", x"1F", x"03", 
															x"FF", x"FF", x"7C", x"00", x"00", x"7C", x"FF", x"FF", x"00", x"00", x"FE", x"C6", x"C6", x"FE", x"00", x"00", x"FF", x"FF", x"00", x"04", x"0C", x"18", x"30", x"00", x"00", x"00", x"06", x"06", x"0C", x"18", x"70", x"60", x"FF", x"FF", x"00", x"04", x"04", x"04", x"08", x"08", x"00", x"00", x"06", x"06", x"04", x"04", x"08", x"08", x"08", x"10", x"10", x"00", x"00", x"10", x"10", x"08", x"08", x"10", x"30", x"30", x"30", x"30", x"10", x"08", x"7F", x"3F", x"3F", x"3E", x"1F", x"0F", x"03", x"00", x"00", x"00", x"01", x"03", x"01", x"00", x"00", x"00", x"03", x"0F", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"03", x"0E", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"22", x"65", x"25", x"25", x"25", x"25", x"77", x"72", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"62", x"95", x"15", x"25", x"45", x"85", x"F7", x"F2", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A2", x"A5", x"A5", x"A5", x"F5", x"F5", x"27", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F2", x"85", x"85", x"E5", x"15", x"15", x"F7", x"E2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"62", x"95", x"55", x"65", x"B5", x"95", x"97", x"62", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"50", x"50", x"50", x"50", x"50", x"70", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"E6", x"66", x"66", x"66", x"67", x"F3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5E", x"59", x"59", x"59", x"5E", x"D8", x"98", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"00", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"06", x"06", x"06", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"18", x"3C", x"3C", x"3C", x"18", x"18", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"7F", x"7F", x"7F", x"FF", x"E3", x"C1", x"FF", x"80", x"80", x"80", x"80", x"00", x"1C", x"3E", x"80", x"80", x"80", x"C1", x"E3", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"3E", x"1C", x"00", x"00", x"FF", x"38", x"7C", x"7C", x"7C", x"7C", x"7C", x"38", x"00", x"08", x"04", x"04", x"04", x"04", x"04", x"08", x"00", x"03", x"06", x"0C", x"0C", x"08", x"08", x"04", x"03", x"03", x"05", x"0B", x"0B", x"0F", x"0F", x"07", x"03", 
															x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"07", x"38", x"C0", x"00", x"00", x"00", x"00", x"00", x"07", x"3F", x"FF", x"00", x"00", x"00", x"00", x"00", x"E0", x"1C", x"03", x"00", x"00", x"00", x"00", x"00", x"E0", x"FC", x"FF", x"80", x"40", x"20", x"10", x"08", x"04", x"02", x"01", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"04", x"0E", x"0E", x"0E", x"6E", x"64", x"60", x"60", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"0F", x"1F", x"1F", x"7F", x"FF", x"FF", x"7F", x"07", x"08", x"10", x"00", x"60", x"80", x"80", x"40", x"03", x"07", x"1F", x"3F", x"3F", x"3F", x"79", x"F7", x"03", x"04", x"18", x"20", x"20", x"20", x"46", x"88", x"C0", x"E0", x"F0", x"F4", x"FE", x"BF", x"DF", x"FF", x"C0", x"20", x"10", x"14", x"0A", x"41", x"21", x"01", 
															x"90", x"B8", x"F8", x"FA", x"FF", x"FF", x"FF", x"FE", x"90", x"A8", x"48", x"0A", x"05", x"01", x"01", x"02", x"3B", x"1D", x"0E", x"0F", x"07", x"00", x"00", x"00", x"24", x"12", x"09", x"08", x"07", x"00", x"00", x"00", x"FF", x"BF", x"1C", x"C0", x"F3", x"FF", x"7E", x"1C", x"00", x"40", x"E3", x"3F", x"0C", x"81", x"62", x"1C", x"BF", x"7F", x"3D", x"83", x"C7", x"FF", x"FF", x"3C", x"40", x"80", x"C2", x"7C", x"38", x"00", x"C3", x"3C", x"FC", x"FE", x"FF", x"FE", x"FE", x"F8", x"60", x"00", x"04", x"02", x"01", x"00", x"06", x"98", x"60", x"00", x"C0", x"20", x"10", x"10", x"10", x"10", x"20", x"C0", x"C0", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"3F", x"7F", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"88", x"9C", x"88", x"80", x"80", x"80", x"80", x"80", x"7F", x"7F", x"7F", x"3E", x"1C", x"00", x"00", x"00", 
															x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"08", x"14", x"24", x"C4", x"03", x"40", x"A1", x"26", x"00", x"08", x"18", x"38", x"FC", x"BF", x"5E", x"D9", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"7F", x"80", x"80", x"98", x"9C", x"8C", x"80", x"80", x"00", x"7F", x"7F", x"67", x"67", x"7F", x"7F", x"7F", x"FF", x"01", x"01", x"FF", x"10", x"10", x"10", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"01", x"01", x"01", x"FF", x"10", x"10", x"10", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"01", x"01", x"19", x"1D", x"0D", x"01", x"01", x"00", x"FF", x"FF", x"E7", x"E7", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"60", x"40", x"C0", x"80", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"80", x"80", x"80", x"80", x"80", x"81", x"42", x"3C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"7C", x"00", x"00", x"00", x"00", x"00", x"01", x"82", x"7C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"7C", x"00", x"00", x"00", x"00", x"00", x"01", x"83", x"FF", 
															x"F8", x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"F8", x"04", x"02", x"02", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"01", x"01", x"01", x"01", x"01", x"81", x"42", x"3C", x"00", x"08", x"08", x"08", x"10", x"10", x"10", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7F", x"7F", x"78", x"73", x"73", x"73", x"7F", x"7F", x"80", x"A0", x"87", x"8F", x"8E", x"8E", x"86", x"00", x"FF", x"FF", x"3F", x"9F", x"9F", x"9F", x"1F", x"FE", x"01", x"05", x"C1", x"E1", x"71", x"71", x"F1", x"7E", x"7E", x"7F", x"7E", x"7E", x"7F", x"7F", x"FF", x"81", x"81", x"80", x"81", x"81", x"A0", x"80", x"FF", x"7F", x"7F", x"FF", x"7F", x"7F", x"FF", x"FF", x"FF", x"F1", x"C1", x"C1", x"81", x"C1", x"C5", x"01", x"FF", x"7F", x"80", x"A0", x"80", x"80", x"80", x"80", x"80", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FE", x"01", x"05", x"01", x"01", x"01", x"01", x"01", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"A0", x"80", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"01", x"01", x"01", x"01", x"01", x"05", x"01", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"FC", x"FE", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"7C", x"11", x"39", x"11", x"01", x"01", x"01", x"01", x"01", x"FE", x"FE", x"FE", x"7C", x"38", x"00", x"00", x"00", x"EF", x"28", x"28", x"28", x"28", x"28", x"EF", x"00", x"20", x"E7", x"E7", x"E7", x"E7", x"E7", x"EF", x"00", x"FE", x"82", x"82", x"82", x"82", x"82", x"FE", x"00", x"02", x"7E", x"7E", x"7E", x"7E", x"7E", x"FE", x"00", x"80", x"80", x"80", x"98", x"9C", x"8C", x"80", x"7F", x"7F", x"7F", x"7F", x"67", x"67", x"7F", x"7F", x"7F", 
															x"FF", x"FF", x"83", x"F3", x"F3", x"F3", x"F3", x"F3", x"FF", x"80", x"FC", x"8C", x"8C", x"8C", x"8C", x"8C", x"FF", x"FF", x"F0", x"F6", x"F6", x"F6", x"F6", x"F6", x"FF", x"00", x"0F", x"09", x"09", x"09", x"09", x"09", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"57", x"2F", x"57", x"2F", x"57", x"FF", x"01", x"FF", x"A9", x"D1", x"A9", x"D1", x"A9", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"FF", x"3F", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"FF", x"3F", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"FF", x"FF", x"09", x"09", x"09", x"09", x"09", x"09", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"2F", x"57", x"2F", x"57", x"2F", x"57", x"FF", x"FC", x"D1", x"A9", x"D1", x"A9", x"D1", x"A9", x"FF", x"FC", 
															x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"23", x"23", x"23", x"23", x"23", x"23", x"23", x"23", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"BC", x"5C", x"BC", x"5C", x"BC", x"5C", x"BC", x"5C", x"44", x"A4", x"44", x"A4", x"44", x"A4", x"44", x"A4", x"1F", x"20", x"40", x"40", x"80", x"80", x"80", x"81", x"1F", x"3F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FE", x"FF", x"80", x"80", x"C0", x"FF", x"FF", x"FE", x"FE", x"FF", x"7F", x"7F", x"3F", x"00", x"00", x"01", x"01", x"FF", x"7F", x"7F", x"FF", x"FF", x"07", x"03", x"03", x"FF", x"80", x"80", x"00", x"00", x"F8", x"FC", x"FC", x"FF", x"00", x"00", x"00", x"00", x"81", x"C3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"3C", x"00", x"F8", x"FC", x"FE", x"FE", x"E3", x"C1", x"81", x"81", x"F8", x"04", x"02", x"02", x"1D", x"3F", x"7F", x"7F", 
															x"83", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"1F", x"FC", x"80", x"80", x"80", x"80", x"80", x"60", x"1F", x"FC", x"FC", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"03", x"03", x"03", x"03", x"01", x"01", x"00", x"FF", x"01", x"01", x"01", x"01", x"03", x"03", x"07", x"FF", x"FE", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"81", x"C1", x"E3", x"FF", x"FF", x"FF", x"FF", x"FE", x"7F", x"3F", x"1D", x"01", x"01", x"01", x"03", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"B5", x"CE", x"80", x"80", x"80", x"80", x"80", x"84", x"CA", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"AD", x"73", x"01", x"01", x"01", x"01", x"01", x"21", x"53", x"8D", x"77", x"77", x"77", x"77", x"77", x"77", x"77", x"77", x"00", x"00", x"00", x"00", x"77", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"77", x"77", x"77", x"77", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"77", x"77", x"77", x"77", x"77", x"01", x"01", x"01", x"19", x"1D", x"0D", x"01", x"FE", x"FF", x"FF", x"FF", x"E7", x"E7", x"FF", x"FF", x"FE", x"20", x"78", x"7F", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"21", x"21", x"41", x"41", x"41", x"41", x"41", x"04", x"9A", x"FA", x"FD", x"FD", x"FD", x"FD", x"FD", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7E", x"38", x"21", x"00", x"01", x"00", x"01", x"00", x"21", x"21", x"01", x"01", x"01", x"01", x"01", x"01", x"FA", x"8A", x"84", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"02", x"04", x"00", x"10", x"00", x"40", x"80", x"00", x"01", x"01", x"06", x"08", x"18", x"20", x"20", x"C0", 
															x"0B", x"0B", x"3B", x"0B", x"FB", x"0B", x"0B", x"0A", x"04", x"04", x"C4", x"F4", x"F4", x"04", x"04", x"05", x"90", x"10", x"1F", x"10", x"1F", x"10", x"10", x"90", x"70", x"F0", x"F0", x"FF", x"FF", x"F0", x"F0", x"70", x"3F", x"78", x"E7", x"CF", x"58", x"58", x"50", x"90", x"C0", x"87", x"18", x"B0", x"E7", x"E7", x"EF", x"EF", x"B0", x"FC", x"E2", x"C1", x"C1", x"83", x"8F", x"7E", x"6F", x"43", x"5D", x"3F", x"3F", x"7F", x"7F", x"FF", x"FE", x"03", x"0F", x"91", x"70", x"60", x"20", x"31", x"03", x"FF", x"F1", x"6E", x"CF", x"DF", x"FF", x"FF", x"3F", x"3F", x"1D", x"39", x"7B", x"F3", x"86", x"FE", x"FD", x"FB", x"FB", x"F7", x"F7", x"0F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"FF", x"FF", x"80", x"80", x"80", x"80", x"FF", x"FF", x"80", x"FE", x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"FF", x"FE", x"03", x"03", x"03", x"03", x"FF", x"FF", x"03", 
															x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"3C", x"FC", x"FC", x"FC", x"FC", x"FC", x"04", x"04", x"23", x"F3", x"0B", x"0B", x"0B", x"07", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"FF", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"03", x"FF", x"FF", x"FF", x"03", x"03", x"03", x"03", x"FF", x"03", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FC", x"FC", x"FE", x"FE", x"FE", x"02", x"FE", x"FE", x"07", x"07", x"03", x"03", x"03", x"FF", x"03", x"03", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"02", x"02", x"02", x"02", x"02", x"02", x"04", x"04", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"AA", x"D5", x"AA", x"FF", x"FF", x"FF", x"FF", x"FF", x"D5", x"AA", x"D5", x"80", x"80", x"FF", x"03", x"03", x"AB", x"57", x"AB", x"FF", x"FF", x"FE", x"FF", x"FF", x"57", x"AB", x"57", x"03", x"03", x"FE", x"00", x"55", x"AA", x"55", x"FF", x"FF", x"FF", x"00", x"FF", x"AA", x"55", x"AA", x"00", x"00", x"FF", x"00", x"04", x"54", x"AC", x"5C", x"FC", x"FC", x"FC", x"3C", x"FF", x"AF", x"57", x"AB", x"0B", x"0B", x"F3", x"23", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"7C", x"7C", x"78", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FE", x"FC", x"FC", x"F8", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"3F", x"FF", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E1", x"F9", x"FD", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"00", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"1F", x"10", x"10", x"10", x"10", x"10", x"10", x"FF", x"00", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"92", x"92", x"92", x"FE", x"FE", x"00", x"00", x"00", x"48", x"48", x"6C", x"00", x"00", x"00", x"FE", x"00", 
															x"0A", x"0A", x"3A", x"0A", x"FB", x"0B", x"0B", x"0B", x"05", x"05", x"C5", x"F5", x"F4", x"04", x"04", x"04", x"90", x"90", x"9F", x"90", x"9F", x"90", x"90", x"90", x"70", x"70", x"70", x"7F", x"7F", x"70", x"70", x"70", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"88", x"91", x"D1", x"53", x"53", x"73", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"BE", x"CE", x"00", x"00", x"07", x"0F", x"0C", x"1B", x"1B", x"1B", x"00", x"00", x"00", x"00", x"03", x"04", x"04", x"04", x"00", x"00", x"E0", x"F0", x"F0", x"F8", x"F8", x"F8", x"00", x"00", x"60", x"30", x"30", x"98", x"98", x"98", x"1B", x"1B", x"1B", x"1B", x"1B", x"0F", x"0F", x"07", x"04", x"04", x"04", x"04", x"04", x"03", x"00", x"00", 
															x"F8", x"F8", x"F8", x"F8", x"F8", x"F0", x"F0", x"E0", x"98", x"98", x"98", x"98", x"98", x"30", x"30", x"60", x"F1", x"11", x"11", x"1F", x"10", x"10", x"10", x"FF", x"0F", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"E0", x"1F", x"10", x"10", x"F0", x"10", x"10", x"10", x"FF", x"E0", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"0F", x"7F", x"BF", x"DF", x"EF", x"F0", x"F0", x"F0", x"F0", x"80", x"40", x"20", x"10", x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F", x"1F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F", x"01", x"03", x"07", x"0F", x"FF", x"FF", x"FF", x"FF", x"0F", x"0F", x"0F", x"0F", x"F7", x"FB", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"1F", x"3F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"1F", x"20", x"40", x"40", x"40", x"80", x"82", x"82", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"3F", x"1E", x"82", x"80", x"A0", x"44", x"43", x"40", x"21", x"1E", x"F8", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"F8", x"04", x"02", x"02", x"02", x"01", x"41", x"41", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FC", x"78", x"41", x"01", x"05", x"22", x"C2", x"02", x"84", x"78", x"7F", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"DE", x"61", x"61", x"61", x"71", x"5E", x"7F", x"61", x"61", x"DF", x"DF", x"DF", x"DF", x"FF", x"C1", x"DF", x"80", x"80", x"C0", x"F0", x"BF", x"8F", x"81", x"7E", x"7F", x"7F", x"FF", x"3F", x"4F", x"71", x"7F", x"FF", x"61", x"61", x"C1", x"C1", x"81", x"81", x"83", x"FE", x"DF", x"DF", x"BF", x"BF", x"7F", x"7F", x"7F", x"7F", 
															x"00", x"00", x"03", x"0F", x"1F", x"3F", x"7F", x"7F", x"00", x"00", x"03", x"0C", x"10", x"20", x"40", x"40", x"00", x"00", x"C0", x"F0", x"F8", x"FC", x"FE", x"FE", x"00", x"00", x"C0", x"30", x"08", x"04", x"02", x"02", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"7F", x"7F", x"7F", x"3F", x"3F", x"1F", x"0F", x"07", x"40", x"40", x"40", x"20", x"30", x"1C", x"0F", x"07", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"F0", x"F0", x"02", x"02", x"02", x"04", x"0C", x"38", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"07", x"0F", x"08", x"08", x"08", x"08", x"08", x"0C", x"05", x"0A", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"F0", x"10", x"50", x"50", x"50", x"50", x"30", x"A0", x"50", 
															x"81", x"C1", x"A3", x"A3", x"9D", x"81", x"81", x"81", x"00", x"41", x"22", x"22", x"1C", x"00", x"00", x"00", x"E3", x"F7", x"C1", x"C1", x"C1", x"C1", x"F7", x"E3", x"E3", x"14", x"3E", x"3E", x"3E", x"3E", x"14", x"E3", x"00", x"00", x"07", x"0F", x"0C", x"1B", x"1B", x"1B", x"FF", x"FF", x"F8", x"F0", x"F0", x"E0", x"E0", x"E0", x"00", x"00", x"E0", x"F0", x"F0", x"F8", x"F8", x"F8", x"FF", x"FF", x"7F", x"3F", x"3F", x"9F", x"9F", x"9F", x"1B", x"1B", x"1B", x"1B", x"1B", x"0F", x"0F", x"07", x"E0", x"E0", x"E0", x"E0", x"E0", x"F3", x"F0", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F0", x"F0", x"E0", x"9F", x"9F", x"9F", x"9F", x"9F", x"3F", x"3F", x"7F", x"E0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"70", x"1F", x"10", x"70", x"7F", x"7F", x"7F", x"07", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"03", x"F8", x"00", x"03", x"FB", x"FB", x"FB", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"EF", x"7C", x"7B", x"76", x"75", x"75", x"77", x"17", x"67", x"FF", x"DF", x"EF", x"AF", x"AF", x"6F", x"EF", x"E7", x"3B", x"FB", x"7B", x"FB", x"FB", x"F3", x"F8", x"F3", x"1F", x"1F", x"3F", x"3F", x"70", x"63", x"E7", x"E5", x"0F", x"0F", x"1F", x"1F", x"3F", x"3C", x"78", x"7A", x"F0", x"F0", x"F8", x"F8", x"0C", x"C4", x"E4", x"A6", x"F8", x"F8", x"FC", x"FC", x"FE", x"3E", x"1E", x"5F", x"E9", x"E9", x"E9", x"EF", x"E2", x"E3", x"F0", x"FF", x"76", x"76", x"76", x"70", x"7D", x"7C", x"7F", x"7F", x"96", x"96", x"96", x"F6", x"46", x"C6", x"0E", x"FE", x"6F", x"6F", x"6F", x"0F", x"BF", x"3F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"3C", x"3C", x"7E", x"7E", x"FF", x"FF", x"FF", x"42", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"0F", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"7F", x"F0", x"E0", x"E0", x"C0", x"C0", x"80", x"80", x"80", x"F0", x"F8", x"F8", x"FC", x"FC", x"FE", x"FE", x"FE", x"0F", x"07", x"07", x"03", x"03", x"01", x"01", x"01", x"7F", x"7F", x"3F", x"3F", x"3F", x"3F", x"1F", x"1F", x"80", x"80", x"C0", x"C0", x"E0", x"F8", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FC", x"FC", x"FE", x"FE", x"FF", x"7F", x"1F", x"07", x"03", x"03", x"01", x"81", x"7F", x"7F", x"7F", x"3F", x"3F", x"3F", x"3F", x"1F", x"80", x"80", x"80", x"C0", x"C0", x"E0", x"E0", x"F0", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"01", x"01", x"01", x"03", x"03", x"07", x"07", x"0F", x"1F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"FC", x"F8", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"7E", x"7E", x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"01", x"01", x"01", x"03", x"03", x"07", x"07", x"0F", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"FF", x"FF", x"FF", x"FF", x"FC", x"FE", x"FE", x"7E", x"FF", x"03", x"03", x"03", x"03", x"03", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"01", x"01", x"01", x"03", x"07", x"03", x"01", x"01", 
															x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"7C", x"7C", x"78", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"7F", x"7F", x"3F", x"3F", x"3F", x"3F", x"1F", x"1F", x"80", x"80", x"C0", x"C0", x"E0", x"F8", x"FE", x"FF", x"3F", x"BF", x"FF", x"FF", x"FC", x"FC", x"FE", x"FE", x"FF", x"7F", x"1F", x"07", x"03", x"03", x"01", x"81", x"7F", x"7F", x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"7E", x"7E", x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"81", x"81", x"81", x"81", x"81", x"81", x"81", x"81", 
															x"81", x"C3", x"C3", x"E7", x"E7", x"FF", x"FF", x"FF", x"7E", x"3C", x"3C", x"18", x"18", x"00", x"00", x"00", x"0F", x"43", x"5B", x"53", x"31", x"19", x"0F", x"07", x"F2", x"FE", x"FE", x"FF", x"FF", x"EF", x"F7", x"F8", x"C1", x"C3", x"C6", x"84", x"FC", x"FC", x"0E", x"02", x"BF", x"BE", x"BD", x"7B", x"7B", x"07", x"F3", x"FD", x"10", x"20", x"22", x"BA", x"E6", x"E1", x"C0", x"C0", x"FF", x"FF", x"FF", x"67", x"59", x"9E", x"BF", x"BF", x"20", x"A6", x"54", x"26", x"20", x"C6", x"54", x"26", x"20", x"E6", x"54", x"26", x"21", x"06", x"54", x"26", x"20", x"85", x"01", x"44", x"20", x"86", x"54", x"48", x"20", x"9A", x"01", x"49", x"20", x"A5", x"C9", x"46", x"20", x"BA", x"C9", x"4A", x"20", x"A6", x"0A", x"D0", x"D1", x"D8", x"D8", x"DE", x"D1", x"D0", x"DA", x"DE", x"D1", x"20", x"C6", x"0A", x"D2", x"D3", x"DB", x"DB", x"DB", x"D9", x"DB", x"DC", x"DB", x"DF", x"20", x"E6", 
															x"0A", x"D4", x"D5", x"D4", x"D9", x"DB", x"E2", x"D4", x"DA", x"DB", x"E0", x"21", x"06", x"0A", x"D6", x"D7", x"D6", x"D7", x"E1", x"26", x"D6", x"DD", x"E1", x"E1", x"21", x"26", x"14", x"D0", x"E8", x"D1", x"D0", x"D1", x"DE", x"D1", x"D8", x"D0", x"D1", x"26", x"DE", x"D1", x"DE", x"D1", x"D0", x"D1", x"D0", x"D1", x"26", x"21", x"46", x"14", x"DB", x"42", x"42", x"DB", x"42", x"DB", x"42", x"DB", x"DB", x"42", x"26", x"DB", x"42", x"DB", x"42", x"DB", x"42", x"DB", x"42", x"26", x"21", x"66", x"46", x"DB", x"21", x"6C", x"0E", x"DF", x"DB", x"DB", x"DB", x"26", x"DB", x"DF", x"DB", x"DF", x"DB", x"DB", x"E4", x"E5", x"26", x"21", x"86", x"14", x"DB", x"DB", x"DB", x"DE", x"43", x"DB", x"E0", x"DB", x"DB", x"DB", x"26", x"DB", x"E3", x"DB", x"E0", x"DB", x"DB", x"E6", x"E3", x"26", x"21", x"A6", x"14", x"DB", x"DB", x"DB", x"DB", x"42", x"DB", x"DB", x"DB", x"D4", x"D9", x"26", 
															x"DB", x"D9", x"DB", x"DB", x"D4", x"D9", x"D4", x"D9", x"E7", x"21", x"C5", x"16", x"5F", x"95", x"95", x"95", x"95", x"95", x"95", x"95", x"95", x"97", x"98", x"78", x"95", x"96", x"95", x"95", x"97", x"98", x"97", x"98", x"95", x"7A", x"21", x"ED", x"0E", x"CF", x"01", x"09", x"08", x"05", x"24", x"17", x"12", x"17", x"1D", x"0E", x"17", x"0D", x"18", x"22", x"4B", x"0D", x"01", x"24", x"19", x"15", x"0A", x"22", x"0E", x"1B", x"24", x"10", x"0A", x"16", x"0E", x"22", x"8B", x"0D", x"02", x"24", x"19", x"15", x"0A", x"22", x"0E", x"1B", x"24", x"10", x"0A", x"16", x"0E", x"22", x"EC", x"04", x"1D", x"18", x"19", x"28", x"22", x"F6", x"01", x"00", x"23", x"C9", x"56", x"55", x"23", x"E2", x"04", x"99", x"AA", x"AA", x"AA", x"23", x"EA", x"04", x"99", x"AA", x"AA", x"AA", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF");
	
	type AUDIO_TEST_ARRAY is array (0 to 9399) of unsigned(7 downto 0);
	constant AUDIO_ROM : AUDIO_TEST_ARRAY := (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FD",x"FD",x"FE",x"FE",x"FC",x"FC",x"FF",x"05",x"0C",x"0F",x"0C",x"04",x"F9",x"EF",x"E9",x"EC",x"F8",x"07",x"14",x"1B",x"1A",x"0D",x"FA",x"E7",x"D8",x"D1",x"D6",x"E3",x"F3",x"02",x"0B",x"0A",x"00",x"F4",x"EA",x"E7",x"ED",x"FC",x"0E",x"20",x"2B",x"2D",x"25",x"15",x"03",x"F3",x"E9",x"E9",
															x"F1",x"FA",x"00",x"FF",x"F5",x"E3",x"CE",x"BA",x"AD",x"AB",x"B5",x"C6",x"D9",x"EB",x"F6",x"F7",x"F1",x"E9",x"E7",x"EB",x"F9",x"10",x"29",x"3E",x"4C",x"50",x"49",x"3A",x"29",x"1A",x"13",x"14",x"1D",x"25",x"29",x"24",x"15",x"FD",x"E2",x"CC",x"BE",x"BD",x"C7",x"D8",x"EA",x"F9",x"FF",x"FB",x"F1",x"E8",x"E5",x"EB",x"FB",x"13",x"2B",x"3F",x"4A",x"4B",x"3F",x"2C",x"19",x"0B",x"04",x"05",x"0D",x"16",x"1B",x"17",x"0A",x"F4",x"DB",x"C4",x"B6",x"B2",x"B9",x"C7",x"D9",x"EA",x"F4",x"F5",x"EF",x"E7",x"E4",x"E7",x"F5",x"0B",x"25",x"3B",x"49",x"4B",x"42",x"32",x"21",x"13",x"0B",x"0D",x"14",x"1B",x"1D",x"17",
															x"06",x"EF",x"D6",x"C2",x"B7",x"B7",x"C2",x"D2",x"E3",x"F0",x"F5",x"F2",x"EA",x"E3",x"E2",x"EA",x"FE",x"18",x"31",x"44",x"4E",x"4C",x"41",x"31",x"20",x"13",x"0C",x"0F",x"16",x"1E",x"20",x"1A",x"0A",x"F2",x"DA",x"C5",x"B8",x"B7",x"C0",x"CF",x"E0",x"EE",x"F3",x"EF",x"E7",x"E1",x"E1",x"EB",x"FF",x"17",x"2F",x"42",x"4B",x"47",x"3C",x"2D",x"1E",x"13",x"11",x"17",x"1F",x"24",x"22",x"15",x"FF",x"E4",x"CC",x"BB",x"B4",x"B9",x"C6",x"D6",x"E4",x"ED",x"EC",x"E4",x"DD",x"D9",x"DD",x"EC",x"03",x"1B",x"31",x"41",x"45",x"3F",x"33",x"26",x"1A",x"13",x"16",x"1D",x"24",x"26",x"20",x"0F",x"F8",x"E1",x"CD",x"C1",
															x"C1",x"CA",x"D8",x"E6",x"F0",x"F2",x"EC",x"E3",x"DC",x"DC",x"E5",x"FA",x"12",x"2A",x"3B",x"43",x"3F",x"33",x"25",x"18",x"0F",x"0F",x"18",x"22",x"28",x"28",x"1B",x"04",x"EA",x"D4",x"C4",x"BF",x"C6",x"D4",x"E2",x"EF",x"F5",x"F2",x"E8",x"DE",x"D8",x"DA",x"E9",x"01",x"1B",x"31",x"40",x"43",x"3A",x"2D",x"1E",x"12",x"0D",x"11",x"1B",x"24",x"28",x"22",x"10",x"F7",x"DD",x"C8",x"BD",x"BE",x"C9",x"D8",x"E6",x"EF",x"F1",x"E9",x"DE",x"D7",x"D7",x"E2",x"F8",x"12",x"2B",x"3D",x"45",x"41",x"34",x"25",x"17",x"10",x"13",x"1D",x"28",x"2E",x"2C",x"1E",x"08",x"EF",x"D8",x"C7",x"C2",x"C8",x"D4",x"E3",x"EF",x"F4",
															x"F0",x"E6",x"DC",x"D7",x"DB",x"EA",x"01",x"1A",x"30",x"3E",x"40",x"37",x"29",x"19",x"0E",x"0C",x"12",x"1D",x"27",x"2A",x"22",x"10",x"F8",x"DE",x"CA",x"BF",x"C1",x"CC",x"DB",x"E9",x"F3",x"F3",x"EB",x"E1",x"DA",x"DA",x"E5",x"FA",x"14",x"2C",x"3E",x"44",x"3E",x"31",x"23",x"16",x"0F",x"11",x"1A",x"23",x"2A",x"29",x"1C",x"05",x"EB",x"D4",x"C4",x"BE",x"C5",x"D2",x"E0",x"ED",x"F3",x"EF",x"E6",x"DD",x"D8",x"DD",x"EE",x"06",x"1F",x"34",x"40",x"40",x"37",x"29",x"1B",x"10",x"0E",x"14",x"1F",x"28",x"2B",x"23",x"0F",x"F6",x"DC",x"C8",x"BF",x"C2",x"CE",x"DC",x"EB",x"F4",x"F4",x"EE",x"E4",x"DC",x"DD",x"EA",
															x"00",x"17",x"2C",x"3B",x"41",x"3B",x"2F",x"22",x"15",x"0D",x"0E",x"14",x"1E",x"25",x"25",x"19",x"05",x"ED",x"D7",x"C7",x"C2",x"C8",x"D5",x"E3",x"EF",x"F4",x"F1",x"E9",x"E0",x"DB",x"DF",x"EF",x"05",x"1D",x"33",x"3F",x"3F",x"36",x"28",x"1B",x"11",x"0E",x"13",x"1C",x"24",x"28",x"20",x"0D",x"F6",x"DF",x"CD",x"C5",x"C9",x"D5",x"E4",x"F1",x"F8",x"F7",x"EF",x"E5",x"DE",x"DE",x"EA",x"FE",x"15",x"2B",x"3C",x"41",x"3C",x"30",x"22",x"15",x"0F",x"11",x"19",x"22",x"29",x"27",x"1A",x"06",x"EE",x"D9",x"CC",x"CA",x"D2",x"DF",x"ED",x"F6",x"F9",x"F4",x"EB",x"E2",x"DE",x"E3",x"F3",x"08",x"1E",x"30",x"3A",x"38",
															x"2F",x"22",x"16",x"0E",x"0E",x"15",x"1F",x"27",x"29",x"20",x"0E",x"F8",x"E3",x"D4",x"CE",x"D4",x"DF",x"EC",x"F6",x"FB",x"F8",x"F0",x"E7",x"E1",x"E2",x"ED",x"FF",x"15",x"28",x"34",x"37",x"2F",x"23",x"16",x"0D",x"0A",x"0F",x"18",x"21",x"26",x"23",x"15",x"01",x"EC",x"DA",x"D0",x"D1",x"D9",x"E5",x"F0",x"F9",x"FA",x"F4",x"EC",x"E5",x"E2",x"E7",x"F6",x"0A",x"1E",x"2E",x"35",x"32",x"28",x"1C",x"12",x"0C",x"0D",x"14",x"1C",x"22",x"23",x"1A",x"0A",x"F7",x"E4",x"D7",x"D1",x"D5",x"DE",x"E9",x"F3",x"F9",x"F8",x"F1",x"EA",x"E4",x"E4",x"EE",x"FE",x"12",x"23",x"2F",x"32",x"2C",x"22",x"18",x"10",x"0E",x"12",
															x"19",x"20",x"24",x"21",x"15",x"03",x"EF",x"DE",x"D4",x"D3",x"DA",x"E4",x"EE",x"F5",x"F6",x"F2",x"EA",x"E3",x"E1",x"E7",x"F5",x"08",x"1B",x"2A",x"31",x"2F",x"27",x"1E",x"16",x"11",x"11",x"16",x"1C",x"22",x"23",x"1B",x"0D",x"FB",x"E9",x"DA",x"D5",x"D7",x"DF",x"E8",x"F0",x"F5",x"F3",x"EE",x"E8",x"E4",x"E5",x"EE",x"FD",x"0E",x"1E",x"29",x"2C",x"28",x"20",x"18",x"11",x"0F",x"12",x"17",x"1D",x"20",x"1C",x"10",x"00",x"EF",x"E0",x"D8",x"D9",x"DF",x"E8",x"F0",x"F5",x"F5",x"F0",x"EA",x"E5",x"E4",x"EB",x"F8",x"08",x"18",x"24",x"2A",x"29",x"23",x"1A",x"13",x"0F",x"10",x"14",x"1A",x"1E",x"1E",x"16",x"09",
															x"F8",x"E9",x"DE",x"DB",x"DE",x"E5",x"ED",x"F3",x"F4",x"F1",x"EC",x"E7",x"E4",x"E7",x"F1",x"FF",x"0E",x"1C",x"25",x"26",x"22",x"1B",x"14",x"10",x"10",x"14",x"1A",x"1F",x"20",x"1B",x"0F",x"00",x"F1",x"E5",x"DE",x"DF",x"E4",x"EC",x"F2",x"F4",x"F1",x"EB",x"E6",x"E2",x"E2",x"E9",x"F6",x"05",x"14",x"1F",x"24",x"22",x"1C",x"15",x"0F",x"0E",x"11",x"17",x"1C",x"1F",x"1E",x"15",x"08",x"F9",x"EB",x"E2",x"DF",x"E2",x"E9",x"F0",x"F4",x"F4",x"F1",x"EB",x"E5",x"E3",x"E7",x"F1",x"FF",x"0D",x"19",x"21",x"21",x"1C",x"15",x"0F",x"0B",x"0D",x"12",x"18",x"1C",x"1D",x"18",x"0D",x"FF",x"F1",x"E7",x"E2",x"E3",x"E8",
															x"EF",x"F4",x"F7",x"F5",x"F0",x"EB",x"E7",x"E8",x"EE",x"F9",x"07",x"13",x"1C",x"1F",x"1C",x"16",x"10",x"0B",x"0B",x"0E",x"13",x"18",x"1A",x"19",x"11",x"05",x"F9",x"EE",x"E6",x"E5",x"E8",x"EE",x"F4",x"F7",x"F7",x"F3",x"EE",x"EA",x"E8",x"EC",x"F5",x"01",x"0D",x"16",x"1B",x"1B",x"16",x"11",x"0D",x"0B",x"0D",x"12",x"16",x"19",x"19",x"14",x"0B",x"FF",x"F5",x"EC",x"E8",x"E9",x"EC",x"F1",x"F5",x"F6",x"F4",x"EF",x"EB",x"E9",x"EA",x"F0",x"FA",x"05",x"0F",x"17",x"19",x"17",x"13",x"0F",x"0D",x"0E",x"11",x"14",x"17",x"18",x"16",x"0F",x"05",x"FA",x"F0",x"EA",x"E9",x"EB",x"EF",x"F3",x"F4",x"F3",x"EF",x"EB",
															x"E8",x"E8",x"ED",x"F5",x"00",x"0A",x"13",x"17",x"17",x"14",x"10",x"0D",x"0D",x"0F",x"12",x"16",x"18",x"18",x"14",x"0B",x"01",x"F7",x"EF",x"EC",x"EC",x"EF",x"F3",x"F6",x"F6",x"F3",x"EF",x"EC",x"EA",x"EB",x"F2",x"FB",x"05",x"0E",x"15",x"17",x"15",x"12",x"0E",x"0C",x"0C",x"0F",x"12",x"14",x"15",x"13",x"0C",x"03",x"F9",x"F1",x"EC",x"EB",x"ED",x"F0",x"F3",x"F5",x"F4",x"F1",x"EE",x"EC",x"EC",x"F0",x"F8",x"01",x"09",x"11",x"15",x"15",x"13",x"0F",x"0C",x"0B",x"0C",x"0F",x"12",x"15",x"14",x"10",x"09",x"00",x"F7",x"F0",x"ED",x"EE",x"F1",x"F4",x"F6",x"F6",x"F4",x"F1",x"EE",x"EC",x"EE",x"F3",x"FB",x"04",
															x"0C",x"11",x"13",x"11",x"0E",x"0A",x"08",x"09",x"0C",x"10",x"13",x"14",x"12",x"0C",x"04",x"FB",x"F4",x"F0",x"F0",x"F2",x"F6",x"F9",x"FA",x"F8",x"F5",x"F1",x"EF",x"EE",x"F2",x"F8",x"00",x"09",x"0F",x"11",x"11",x"0E",x"0A",x"07",x"07",x"09",x"0D",x"10",x"13",x"12",x"0D",x"06",x"FE",x"F6",x"F1",x"EF",x"F1",x"F4",x"F7",x"FA",x"F9",x"F6",x"F3",x"F1",x"F0",x"F1",x"F7",x"FE",x"06",x"0D",x"10",x"11",x"0E",x"0B",x"08",x"07",x"09",x"0C",x"0F",x"11",x"11",x"0E",x"08",x"01",x"F9",x"F4",x"F1",x"F2",x"F4",x"F7",x"FA",x"FB",x"F9",x"F6",x"F2",x"F0",x"F0",x"F3",x"F9",x"00",x"07",x"0C",x"0E",x"0D",x"0A",x"07",
															x"05",x"06",x"08",x"0B",x"0E",x"10",x"0F",x"0B",x"05",x"FE",x"F8",x"F4",x"F3",x"F5",x"F8",x"FA",x"FC",x"FA",x"F7",x"F4",x"F1",x"F0",x"F2",x"F7",x"FD",x"04",x"0A",x"0D",x"0D",x"0B",x"08",x"05",x"05",x"07",x"0A",x"0D",x"0F",x"10",x"0D",x"08",x"01",x"FB",x"F6",x"F4",x"F4",x"F7",x"FA",x"FC",x"FC",x"F9",x"F6",x"F3",x"F1",x"F2",x"F5",x"FA",x"01",x"07",x"0B",x"0D",x"0C",x"09",x"07",x"05",x"05",x"08",x"0B",x"0E",x"0F",x"0E",x"0A",x"04",x"FE",x"F9",x"F5",x"F4",x"F5",x"F7",x"FA",x"FB",x"FA",x"F7",x"F4",x"F2",x"F1",x"F3",x"F8",x"FD",x"03",x"08",x"0B",x"0C",x"0A",x"08",x"06",x"05",x"07",x"0A",x"0C",x"0E",
															x"0F",x"0D",x"08",x"02",x"FD",x"F8",x"F5",x"F5",x"F6",x"F9",x"FA",x"FA",x"F9",x"F6",x"F3",x"F2",x"F2",x"F5",x"FA",x"FF",x"05",x"09",x"0B",x"0A",x"08",x"06",x"04",x"05",x"08",x"0B",x"0D",x"0F",x"0E",x"0A",x"05",x"00",x"FB",x"F8",x"F7",x"F8",x"F9",x"FB",x"FB",x"FA",x"F7",x"F5",x"F3",x"F2",x"F4",x"F8",x"FC",x"02",x"06",x"08",x"08",x"07",x"05",x"04",x"04",x"06",x"09",x"0C",x"0D",x"0D",x"0B",x"07",x"02",x"FD",x"F9",x"F8",x"F8",x"F9",x"FB",x"FC",x"FB",x"F9",x"F6",x"F4",x"F3",x"F4",x"F7",x"FC",x"00",x"05",x"08",x"08",x"08",x"06",x"05",x"04",x"06",x"08",x"0B",x"0D",x"0D",x"0C",x"08",x"03",x"FE",x"FA",
															x"F8",x"F8",x"F9",x"FA",x"FC",x"FC",x"FA",x"F7",x"F5",x"F3",x"F3",x"F5",x"F9",x"FE",x"03",x"06",x"08",x"08",x"07",x"05",x"04",x"05",x"07",x"0A",x"0C",x"0D",x"0D",x"0A",x"06",x"01",x"FD",x"FA",x"F8",x"F9",x"FA",x"FC",x"FC",x"FB",x"F9",x"F6",x"F4",x"F3",x"F4",x"F7",x"FB",x"00",x"04",x"07",x"08",x"07",x"06",x"04",x"04",x"06",x"08",x"0B",x"0C",x"0D",x"0B",x"08",x"03",x"FF",x"FB",x"F9",x"F9",x"FA",x"FB",x"FC",x"FC",x"FA",x"F8",x"F5",x"F4",x"F4",x"F6",x"F9",x"FD",x"02",x"05",x"07",x"07",x"06",x"05",x"04",x"04",x"06",x"09",x"0B",x"0C",x"0C",x"09",x"05",x"01",x"FD",x"FA",x"F9",x"F9",x"FA",x"FC",x"FC",
															x"FB",x"F9",x"F7",x"F5",x"F4",x"F6",x"F9",x"FC",x"00",x"04",x"06",x"07",x"06",x"05",x"04",x"04",x"05",x"07",x"0A",x"0B",x"0B",x"09",x"06",x"02",x"FF",x"FB",x"FA",x"FA",x"FB",x"FC",x"FD",x"FC",x"FB",x"F8",x"F6",x"F5",x"F5",x"F8",x"FB",x"FF",x"03",x"05",x"06",x"06",x"05",x"04",x"03",x"04",x"06",x"08",x"0A",x"0B",x"0A",x"07",x"04",x"00",x"FD",x"FB",x"FA",x"FB",x"FC",x"FD",x"FD",x"FC",x"FA",x"F7",x"F5",x"F5",x"F6",x"F9",x"FD",x"01",x"05",x"07",x"07",x"06",x"04",x"03",x"04",x"05",x"08",x"09",x"0A",x"0A",x"08",x"05",x"02",x"FE",x"FC",x"FB",x"FB",x"FC",x"FC",x"FD",x"FC",x"FB",x"F9",x"F7",x"F6",x"F7",
															x"F9",x"FC",x"00",x"03",x"05",x"06",x"05",x"05",x"04",x"04",x"04",x"05",x"07",x"08",x"09",x"09",x"06",x"03",x"00",x"FE",x"FD",x"FC",x"FC",x"FC",x"FC",x"FB",x"FB",x"F9",x"F4",x"F3",x"F5",x"F6",x"F5",x"F5",x"F9",x"03",x"11",x"1C",x"1D",x"16",x"08",x"F8",x"EE",x"ED",x"F3",x"FE",x"07",x"0A",x"04",x"F8",x"E9",x"E0",x"DF",x"E6",x"F4",x"04",x"0F",x"10",x"08",x"FA",x"ED",x"E7",x"EA",x"F5",x"06",x"14",x"18",x"12",x"04",x"F3",x"E6",x"E2",x"E7",x"F3",x"00",x"07",x"04",x"F9",x"E9",x"D9",x"D2",x"D4",x"E0",x"EF",x"FC",x"FF",x"F9",x"EB",x"DC",x"D1",x"D0",x"D7",x"E5",x"F7",x"04",x"07",x"01",x"F5",x"E6",x"DE",
															x"DF",x"EA",x"FC",x"0C",x"13",x"11",x"06",x"F6",x"EA",x"E8",x"F0",x"FF",x"11",x"1D",x"1D",x"14",x"03",x"F3",x"EC",x"F0",x"FC",x"0D",x"1B",x"20",x"1A",x"0C",x"FB",x"F0",x"EF",x"F6",x"04",x"13",x"1B",x"19",x"0F",x"FF",x"F1",x"EB",x"EF",x"FC",x"0C",x"17",x"19",x"11",x"04",x"F5",x"EB",x"EA",x"F1",x"FE",x"0E",x"18",x"18",x"0F",x"FF",x"EF",x"E8",x"E9",x"F4",x"05",x"12",x"16",x"10",x"02",x"F1",x"E7",x"E6",x"EF",x"00",x"10",x"17",x"14",x"08",x"F7",x"E9",x"E6",x"EC",x"FB",x"0C",x"16",x"17",x"0E",x"FF",x"F0",x"EA",x"ED",x"F9",x"0A",x"16",x"1A",x"13",x"04",x"F4",x"EB",x"EB",x"F5",x"06",x"14",x"1A",x"16",
															x"0A",x"FB",x"EF",x"EB",x"F0",x"FD",x"0D",x"17",x"18",x"11",x"02",x"F2",x"EA",x"EC",x"F6",x"06",x"13",x"18",x"13",x"06",x"F5",x"EA",x"E9",x"F1",x"00",x"0F",x"18",x"16",x"0B",x"FA",x"EC",x"E6",x"EB",x"F9",x"0B",x"17",x"18",x"10",x"00",x"F0",x"E8",x"EA",x"F5",x"06",x"14",x"18",x"13",x"05",x"F4",x"E8",x"E7",x"F0",x"00",x"11",x"19",x"16",x"0A",x"FA",x"EC",x"E7",x"EC",x"FA",x"0B",x"17",x"19",x"11",x"02",x"F1",x"E9",x"EA",x"F5",x"05",x"14",x"1A",x"15",x"07",x"F6",x"EB",x"E9",x"F1",x"01",x"11",x"1A",x"18",x"0D",x"FC",x"ED",x"E8",x"ED",x"FA",x"0C",x"18",x"19",x"11",x"01",x"F1",x"E8",x"EA",x"F5",x"06",
															x"14",x"19",x"14",x"06",x"F5",x"E9",x"E8",x"F0",x"00",x"11",x"1A",x"18",x"0C",x"FB",x"ED",x"E7",x"EC",x"F9",x"0B",x"17",x"1A",x"12",x"02",x"F1",x"E7",x"E7",x"F2",x"04",x"13",x"1A",x"16",x"08",x"F6",x"E9",x"E7",x"EF",x"FF",x"10",x"1A",x"19",x"0D",x"FC",x"EC",x"E6",x"EB",x"F9",x"0B",x"18",x"1A",x"12",x"02",x"F1",x"E7",x"E9",x"F4",x"05",x"14",x"1A",x"14",x"06",x"F5",x"E9",x"E7",x"F0",x"01",x"12",x"1B",x"18",x"0C",x"FB",x"ED",x"E7",x"EC",x"FA",x"0B",x"18",x"1A",x"12",x"03",x"F2",x"E8",x"E9",x"F4",x"04",x"13",x"1A",x"15",x"09",x"F8",x"EC",x"E9",x"F0",x"FF",x"0F",x"18",x"18",x"0E",x"FE",x"EE",x"E8",
															x"EB",x"F8",x"09",x"16",x"19",x"12",x"03",x"F3",x"EA",x"EA",x"F4",x"03",x"11",x"17",x"13",x"07",x"F7",x"EB",x"E9",x"F0",x"FE",x"0F",x"18",x"16",x"0C",x"FD",x"EF",x"E9",x"EC",x"F7",x"07",x"14",x"19",x"13",x"06",x"F6",x"EB",x"EA",x"F2",x"01",x"10",x"17",x"15",x"0A",x"FA",x"ED",x"E9",x"EF",x"FC",x"0D",x"17",x"18",x"10",x"01",x"F2",x"EA",x"EC",x"F6",x"06",x"13",x"17",x"12",x"05",x"F6",x"ED",x"EC",x"F4",x"02",x"10",x"17",x"14",x"09",x"FA",x"EF",x"EC",x"F1",x"FD",x"0C",x"15",x"16",x"0E",x"00",x"F2",x"EB",x"EE",x"F8",x"07",x"14",x"19",x"14",x"07",x"F7",x"EC",x"EA",x"F2",x"00",x"10",x"18",x"16",x"0C",
															x"FC",x"EF",x"EA",x"EF",x"FC",x"0C",x"17",x"19",x"12",x"04",x"F5",x"EC",x"ED",x"F6",x"05",x"13",x"18",x"14",x"08",x"F9",x"EE",x"EB",x"F2",x"01",x"10",x"17",x"16",x"0C",x"FD",x"F0",x"EC",x"F1",x"FE",x"0C",x"17",x"17",x"0D",x"FD",x"F0",x"E8",x"E9",x"F2",x"FF",x"0A",x"13",x"17",x"19",x"17",x"12",x"0C",x"06",x"00",x"FA",x"F6",x"F1",x"ED",x"E9",x"E7",x"E6",x"E7",x"EA",x"EE",x"F3",x"F8",x"FD",x"01",x"05",x"07",x"09",x"0B",x"0D",x"10",x"13",x"16",x"19",x"1A",x"19",x"17",x"13",x"0D",x"07",x"01",x"FA",x"F4",x"EE",x"E8",x"E3",x"DF",x"DB",x"D9",x"D8",x"D7",x"D6",x"D6",x"D6",x"D7",x"D9",x"DC",x"E1",x"E7",
															x"EE",x"F6",x"FF",x"08",x"10",x"17",x"1D",x"23",x"28",x"2B",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2D",x"2C",x"2A",x"26",x"22",x"1B",x"14",x"0C",x"03",x"FA",x"F2",x"EB",x"E5",x"DF",x"DA",x"D7",x"D5",x"D4",x"D4",x"D3",x"D2",x"D1",x"D1",x"D3",x"D6",x"DB",x"E1",x"E9",x"F1",x"FA",x"02",x"0A",x"12",x"18",x"1E",x"24",x"28",x"2A",x"2C",x"2D",x"2D",x"2E",x"2E",x"2D",x"2C",x"28",x"24",x"1E",x"17",x"0F",x"08",x"00",x"F8",x"F2",x"EC",x"E6",x"E1",x"DC",x"D9",x"D7",x"D5",x"D4",x"D2",x"D1",x"D1",x"D2",x"D4",x"D9",x"DE",x"E6",x"EE",x"F6",x"FE",x"07",x"0F",x"16",x"1D",x"24",x"2A",x"2E",x"31",x"33",x"34",x"36",
															x"37",x"38",x"38",x"35",x"31",x"2C",x"25",x"1D",x"14",x"0B",x"01",x"F8",x"EE",x"E5",x"DD",x"D6",x"D0",x"CD",x"CA",x"C8",x"C6",x"C4",x"C3",x"C3",x"C5",x"C9",x"CF",x"D7",x"E0",x"E9",x"F3",x"FE",x"08",x"11",x"1A",x"23",x"2A",x"2F",x"33",x"35",x"37",x"39",x"3A",x"3B",x"3B",x"39",x"35",x"30",x"29",x"21",x"18",x"0E",x"04",x"F9",x"F0",x"E7",x"DF",x"D8",x"D3",x"D0",x"CE",x"CC",x"CB",x"CA",x"C9",x"C9",x"CB",x"CF",x"D4",x"DB",x"E3",x"EC",x"F5",x"FF",x"09",x"12",x"1B",x"22",x"29",x"2E",x"31",x"33",x"35",x"36",x"38",x"39",x"39",x"37",x"34",x"2F",x"29",x"21",x"18",x"0E",x"03",x"F9",x"F0",x"E7",x"DF",x"D7",
															x"D2",x"CE",x"CC",x"CA",x"C8",x"C6",x"C5",x"C5",x"C6",x"CA",x"CF",x"D6",x"DE",x"E7",x"F2",x"FC",x"07",x"11",x"1A",x"23",x"2A",x"30",x"34",x"37",x"39",x"3A",x"3C",x"3D",x"3C",x"3A",x"37",x"31",x"2A",x"21",x"18",x"0E",x"03",x"F8",x"EF",x"E6",x"DE",x"D7",x"D1",x"CE",x"CC",x"CB",x"CA",x"C9",x"C8",x"C9",x"CA",x"CD",x"D2",x"D9",x"E1",x"EA",x"F4",x"FE",x"08",x"11",x"19",x"21",x"28",x"2D",x"31",x"32",x"33",x"34",x"35",x"36",x"36",x"35",x"32",x"2D",x"27",x"20",x"17",x"0E",x"04",x"FB",x"F2",x"EA",x"E2",x"DC",x"D6",x"D3",x"D1",x"CF",x"CE",x"CD",x"CC",x"CC",x"CC",x"CF",x"D3",x"D8",x"DF",x"E7",x"F0",x"FA",
															x"03",x"0C",x"14",x"1C",x"23",x"29",x"2D",x"2F",x"31",x"33",x"35",x"36",x"37",x"37",x"35",x"31",x"2B",x"24",x"1C",x"13",x"0A",x"00",x"F6",x"EE",x"E6",x"DE",x"D7",x"D3",x"D0",x"CE",x"CC",x"C9",x"C7",x"C6",x"C6",x"C8",x"CB",x"D0",x"D6",x"DF",x"E9",x"F4",x"FF",x"09",x"13",x"1C",x"24",x"2B",x"31",x"35",x"37",x"39",x"3A",x"3C",x"3D",x"3C",x"3A",x"37",x"32",x"2B",x"23",x"19",x"0F",x"04",x"FA",x"F0",x"E7",x"DE",x"D7",x"D1",x"CD",x"CB",x"C9",x"C7",x"C5",x"C4",x"C4",x"C5",x"C9",x"CE",x"D5",x"DD",x"E7",x"F1",x"FC",x"06",x"10",x"1A",x"22",x"2A",x"30",x"34",x"37",x"39",x"3B",x"3C",x"3D",x"3D",x"3B",x"38",
															x"33",x"2C",x"24",x"1B",x"12",x"08",x"FE",x"F4",x"EC",x"E3",x"DC",x"D6",x"D2",x"D0",x"CE",x"CD",x"CB",x"CB",x"CB",x"CC",x"CF",x"D3",x"D9",x"E1",x"E9",x"F3",x"FC",x"06",x"0F",x"18",x"1F",x"26",x"2C",x"30",x"32",x"34",x"35",x"36",x"37",x"36",x"35",x"32",x"2D",x"28",x"20",x"18",x"10",x"07",x"FE",x"F6",x"EE",x"E7",x"E1",x"DC",x"D8",x"D5",x"D4",x"D3",x"D2",x"D1",x"D1",x"D2",x"D5",x"D9",x"DE",x"E4",x"EB",x"F3",x"FB",x"03",x"0A",x"11",x"18",x"1E",x"23",x"26",x"28",x"2A",x"2C",x"2D",x"2E",x"2E",x"2D",x"2B",x"28",x"23",x"1D",x"17",x"10",x"09",x"01",x"FA",x"F3",x"ED",x"E7",x"E2",x"DE",x"DC",x"DB",x"DA",
															x"D8",x"D7",x"D7",x"D8",x"DA",x"DD",x"E1",x"E7",x"ED",x"F4",x"FC",x"03",x"0A",x"10",x"16",x"1B",x"1F",x"22",x"24",x"25",x"26",x"27",x"28",x"28",x"28",x"26",x"23",x"1E",x"19",x"13",x"0C",x"05",x"FF",x"F9",x"F3",x"EE",x"E9",x"E5",x"E3",x"E1",x"E0",x"DF",x"DE",x"DD",x"DC",x"DC",x"DE",x"E1",x"E5",x"EA",x"F0",x"F6",x"FC",x"02",x"08",x"0D",x"12",x"17",x"1A",x"1D",x"1F",x"21",x"22",x"23",x"25",x"25",x"25",x"23",x"21",x"1D",x"18",x"13",x"0D",x"07",x"01",x"FC",x"F7",x"F2",x"EE",x"EA",x"E6",x"E4",x"E3",x"E1",x"E0",x"DF",x"DE",x"DE",x"DE",x"E1",x"E4",x"E8",x"ED",x"F3",x"F9",x"FF",x"05",x"0A",x"0F",x"14",
															x"18",x"1C",x"1E",x"20",x"21",x"23",x"24",x"25",x"25",x"24",x"22",x"1E",x"1A",x"15",x"0F",x"09",x"03",x"FD",x"F7",x"F2",x"ED",x"E9",x"E6",x"E3",x"E2",x"E1",x"E0",x"DF",x"DE",x"DE",x"DF",x"E1",x"E4",x"E8",x"ED",x"F3",x"F9",x"FF",x"05",x"0A",x"0F",x"14",x"18",x"1B",x"1D",x"1F",x"20",x"20",x"21",x"22",x"22",x"21",x"1F",x"1C",x"17",x"13",x"0D",x"08",x"02",x"FC",x"F7",x"F2",x"EE",x"EA",x"E7",x"E5",x"E3",x"E3",x"E2",x"E1",x"E1",x"E1",x"E1",x"E3",x"E6",x"EA",x"EE",x"F3",x"F9",x"FE",x"04",x"0A",x"0E",x"13",x"17",x"1A",x"1C",x"1D",x"1E",x"1E",x"1F",x"20",x"20",x"1F",x"1E",x"1B",x"18",x"14",x"0F",x"0A",
															x"04",x"FF",x"FA",x"F5",x"F1",x"ED",x"EA",x"E7",x"E6",x"E5",x"E4",x"E3",x"E2",x"E2",x"E2",x"E3",x"E6",x"E9",x"ED",x"F2",x"F7",x"FC",x"02",x"07",x"0B",x"10",x"14",x"17",x"19",x"1B",x"1C",x"1D",x"1E",x"1F",x"20",x"1F",x"1E",x"1C",x"18",x"14",x"10",x"0B",x"05",x"00",x"FB",x"F6",x"F2",x"EE",x"EB",x"E8",x"E7",x"E5",x"E4",x"E3",x"E3",x"E2",x"E3",x"E4",x"E7",x"EA",x"EE",x"F3",x"F8",x"FD",x"02",x"07",x"0B",x"0F",x"13",x"16",x"18",x"1A",x"1B",x"1C",x"1C",x"1D",x"1D",x"1C",x"1A",x"18",x"15",x"11",x"0D",x"08",x"04",x"FF",x"FA",x"F6",x"F2",x"EF",x"EC",x"E9",x"E8",x"E7",x"E6",x"E6",x"E5",x"E5",x"E6",x"E7",
															x"EA",x"ED",x"F0",x"F4",x"F9",x"FE",x"02",x"07",x"0B",x"0E",x"12",x"14",x"16",x"18",x"18",x"19",x"19",x"19",x"19",x"19",x"18",x"16",x"13",x"0F",x"0C",x"08",x"03",x"FF",x"FB",x"F7",x"F4",x"F1",x"EE",x"EC",x"EB",x"EA",x"EA",x"E9",x"E9",x"E8",x"E9",x"E9",x"EB",x"ED",x"F0",x"F4",x"F7",x"FC",x"00",x"04",x"08",x"0C",x"0F",x"12",x"14",x"15",x"16",x"16",x"17",x"17",x"17",x"17",x"16",x"15",x"13",x"11",x"0E",x"0A",x"07",x"03",x"FF",x"FC",x"F9",x"F6",x"F3",x"F1",x"EF",x"EE",x"ED",x"EC",x"EB",x"EA",x"EA",x"EA",x"EB",x"ED",x"EF",x"F2",x"F6",x"FA",x"FD",x"01",x"05",x"08",x"0B",x"0E",x"10",x"12",x"13",x"14",
															x"15",x"16",x"16",x"17",x"16",x"15",x"13",x"11",x"0E",x"0B",x"07",x"04",x"00",x"FC",x"F9",x"F6",x"F3",x"F0",x"EF",x"EE",x"ED",x"EC",x"EC",x"EC",x"EC",x"ED",x"EE",x"F0",x"F2",x"F5",x"F8",x"FB",x"FE",x"02",x"05",x"07",x"0A",x"0D",x"0F",x"11",x"12",x"13",x"14",x"14",x"14",x"15",x"14",x"13",x"11",x"0E",x"0B",x"09",x"05",x"00",x"FD",x"FB",x"F8",x"F3",x"EE",x"ED",x"F2",x"FB",x"01",x"00",x"F6",x"E8",x"DC",x"DA",x"E2",x"EF",x"FA",x"FE",x"F8",x"EE",x"E7",x"EA",x"F7",x"07",x"14",x"18",x"12",x"08",x"01",x"00",x"09",x"14",x"1C",x"1B",x"12",x"05",x"FA",x"F7",x"FE",x"07",x"0D",x"0A",x"FD",x"ED",x"E1",x"DF",
															x"E6",x"F0",x"F8",x"F6",x"EA",x"DB",x"D1",x"D1",x"DB",x"E7",x"EE",x"EE",x"E6",x"DC",x"D5",x"D6",x"E0",x"EE",x"FB",x"00",x"FB",x"F2",x"E8",x"E6",x"EF",x"FC",x"08",x"0C",x"06",x"FC",x"F3",x"F2",x"FA",x"07",x"12",x"14",x"0D",x"01",x"F7",x"F7",x"00",x"0D",x"16",x"15",x"0C",x"FF",x"F7",x"F9",x"02",x"0C",x"13",x"11",x"07",x"FC",x"F5",x"F7",x"01",x"0C",x"13",x"11",x"07",x"FB",x"F4",x"F7",x"02",x"0D",x"12",x"0E",x"03",x"F9",x"F2",x"F4",x"FE",x"0A",x"12",x"10",x"06",x"F9",x"EE",x"EE",x"F7",x"04",x"0D",x"0C",x"02",x"F6",x"EE",x"F0",x"FA",x"06",x"0D",x"0A",x"00",x"F5",x"F0",x"F4",x"FE",x"09",x"0F",x"0B",
															x"00",x"F5",x"F2",x"F7",x"03",x"0D",x"0F",x"09",x"FD",x"F3",x"F1",x"F8",x"04",x"0E",x"0F",x"07",x"FC",x"F3",x"F3",x"FC",x"08",x"11",x"10",x"07",x"FB",x"F4",x"F5",x"FF",x"0B",x"13",x"11",x"07",x"FA",x"F1",x"F3",x"FD",x"09",x"11",x"0F",x"05",x"F8",x"F2",x"F5",x"00",x"0C",x"12",x"0E",x"02",x"F7",x"F2",x"F7",x"02",x"0D",x"10",x"0A",x"FF",x"F4",x"F0",x"F7",x"03",x"0D",x"0F",x"07",x"FB",x"F1",x"EF",x"F7",x"03",x"0D",x"0E",x"05",x"F9",x"F0",x"F0",x"FA",x"06",x"0F",x"0E",x"04",x"F9",x"F1",x"F3",x"FD",x"08",x"10",x"0E",x"04",x"F8",x"F0",x"F3",x"FD",x"09",x"10",x"0D",x"03",x"F9",x"F3",x"F6",x"01",x"0C",
															x"11",x"0C",x"01",x"F7",x"F2",x"F8",x"03",x"0D",x"11",x"0B",x"00",x"F6",x"F3",x"FA",x"05",x"0E",x"10",x"09",x"FD",x"F4",x"F3",x"FB",x"05",x"0E",x"0E",x"05",x"FA",x"F2",x"F3",x"FC",x"07",x"0E",x"0C",x"03",x"F9",x"F2",x"F5",x"FF",x"0A",x"10",x"0C",x"02",x"F7",x"F1",x"F4",x"FE",x"0A",x"10",x"0D",x"02",x"F7",x"F2",x"F7",x"01",x"0B",x"10",x"0A",x"FF",x"F5",x"F0",x"F6",x"01",x"0B",x"0E",x"07",x"FC",x"F2",x"F1",x"F8",x"03",x"0D",x"0F",x"08",x"FD",x"F4",x"F3",x"FC",x"07",x"10",x"0F",x"06",x"FB",x"F3",x"F3",x"FC",x"07",x"0F",x"0D",x"03",x"F8",x"F1",x"F5",x"FF",x"0A",x"10",x"0D",x"03",x"F8",x"F1",x"F5",
															x"FF",x"0A",x"11",x"0D",x"03",x"F7",x"F1",x"F5",x"00",x"0B",x"10",x"0B",x"00",x"F5",x"F1",x"F7",x"02",x"0C",x"0F",x"08",x"FD",x"F3",x"F1",x"F8",x"04",x"0D",x"0F",x"07",x"FD",x"F4",x"F4",x"FC",x"07",x"10",x"0F",x"06",x"FB",x"F3",x"F5",x"FD",x"08",x"0F",x"0C",x"02",x"F7",x"F1",x"F5",x"FF",x"09",x"0E",x"0A",x"01",x"F7",x"F1",x"F4",x"FE",x"0A",x"10",x"0D",x"03",x"F8",x"F2",x"F5",x"FF",x"0A",x"0F",x"0B",x"00",x"F6",x"F2",x"F7",x"02",x"0C",x"10",x"0A",x"FF",x"F5",x"F3",x"F9",x"04",x"0D",x"0F",x"08",x"FD",x"F4",x"F3",x"FB",x"06",x"0E",x"0E",x"07",x"FC",x"F4",x"F5",x"FE",x"09",x"10",x"0E",x"06",x"FB",
															x"F4",x"F6",x"FF",x"0A",x"10",x"0C",x"03",x"F9",x"F3",x"F7",x"01",x"0C",x"12",x"0E",x"04",x"F9",x"F3",x"F7",x"00",x"0B",x"0F",x"0B",x"01",x"F7",x"F3",x"F9",x"03",x"0D",x"10",x"0A",x"00",x"F7",x"F5",x"FC",x"06",x"0E",x"0F",x"08",x"FE",x"F6",x"F5",x"FC",x"06",x"0E",x"0D",x"05",x"FB",x"F4",x"F6",x"FE",x"08",x"0F",x"0D",x"05",x"FB",x"F5",x"F8",x"01",x"0A",x"10",x"0C",x"03",x"F9",x"F5",x"F8",x"01",x"0B",x"0F",x"0B",x"02",x"F8",x"F4",x"F8",x"02",x"0B",x"0F",x"0A",x"00",x"F7",x"F5",x"FA",x"04",x"0D",x"0E",x"08",x"FF",x"F7",x"F6",x"FD",x"07",x"0E",x"0E",x"07",x"FD",x"F7",x"F7",x"FE",x"07",x"0D",x"0C",
															x"04",x"FA",x"F5",x"F7",x"FF",x"08",x"0D",x"0A",x"02",x"F9",x"F5",x"F9",x"01",x"0A",x"0E",x"0A",x"02",x"FA",x"F6",x"FA",x"03",x"0A",x"0D",x"08",x"00",x"F8",x"F6",x"FA",x"03",x"0B",x"0D",x"09",x"00",x"F9",x"F7",x"FC",x"05",x"0C",x"0D",x"07",x"FE",x"F7",x"F7",x"FD",x"05",x"0B",x"0B",x"05",x"FD",x"F7",x"F8",x"FF",x"07",x"0C",x"0A",x"03",x"FB",x"F7",x"F9",x"00",x"08",x"0C",x"09",x"01",x"FA",x"F7",x"FA",x"02",x"09",x"0C",x"08",x"01",x"FA",x"F8",x"FC",x"03",x"0A",x"0C",x"08",x"00",x"F8",x"F6",x"FB",x"02",x"09",x"0C",x"07",x"00",x"F9",x"F7",x"FC",x"04",x"0A",x"0B",x"06",x"FE",x"F8",x"F7",x"FD",x"05",
															x"0A",x"0A",x"03",x"FC",x"F7",x"F8",x"FF",x"07",x"0B",x"0A",x"03",x"FB",x"F7",x"FA",x"01",x"08",x"0C",x"09",x"01",x"FA",x"F7",x"FA",x"02",x"09",x"0B",x"07",x"FF",x"F9",x"F6",x"FB",x"03",x"09",x"0A",x"06",x"FF",x"F8",x"F7",x"FC",x"03",x"0A",x"0B",x"06",x"FE",x"F8",x"F7",x"FC",x"04",x"0A",x"0A",x"05",x"FD",x"F8",x"F8",x"FE",x"05",x"0A",x"09",x"03",x"FC",x"F8",x"F9",x"FF",x"06",x"0A",x"08",x"02",x"FB",x"F8",x"FA",x"01",x"07",x"0A",x"07",x"01",x"FA",x"F8",x"FB",x"01",x"07",x"09",x"05",x"FF",x"F9",x"F8",x"FC",x"02",x"08",x"09",x"05",x"FF",x"FA",x"F9",x"FE",x"04",x"09",x"0A",x"05",x"FE",x"F9",x"F8",
															x"FD",x"03",x"08",x"08",x"04",x"FE",x"F9",x"FA",x"FE",x"04",x"08",x"08",x"03",x"FD",x"F9",x"FA",x"FF",x"05",x"08",x"06",x"01",x"FB",x"F8",x"FB",x"00",x"06",x"09",x"06",x"01",x"FB",x"F9",x"FC",x"02",x"07",x"09",x"05",x"FF",x"FA",x"F9",x"FC",x"02",x"07",x"08",x"04",x"FE",x"F9",x"F9",x"FE",x"04",x"08",x"08",x"04",x"FE",x"F9",x"F9",x"FD",x"04",x"08",x"08",x"03",x"FD",x"F9",x"FA",x"FF",x"05",x"09",x"08",x"03",x"FD",x"F9",x"FB",x"00",x"06",x"09",x"07",x"01",x"FB",x"F9",x"FB",x"00",x"06",x"08",x"06",x"00",x"FB",x"F9",x"FC",x"02",x"07",x"08",x"05",x"FF",x"FA",x"F9",x"FD",x"03",x"07",x"08",x"03",x"FE",
															x"F9",x"F9",x"FE",x"03",x"07",x"07",x"03",x"FD",x"F9",x"FA",x"FE",x"04",x"08",x"07",x"03",x"FD",x"F9",x"FA",x"FF",x"05",x"08",x"07",x"02",x"FC",x"F9",x"FB",x"00",x"06",x"08",x"06",x"00",x"FB",x"F9",x"FC",x"01",x"05",x"07",x"04",x"FE",x"FA",x"F9",x"FC",x"02",x"06",x"07",x"03",x"FE",x"FA",x"FB",x"FF",x"04",x"08",x"08",x"04",x"FE",x"FB",x"FC",x"00",x"04",x"07",x"06",x"02",x"FD",x"F9",x"FA",x"FF",x"04",x"07",x"06",x"02",x"FD",x"FA",x"FB",x"FF",x"03",x"06",x"04",x"00",x"FB",x"FA",x"FC",x"01",x"06",x"07",x"05",x"00",x"FC",x"FA",x"FD",x"01",x"05",x"06",x"04",x"FF",x"FB",x"FA",x"FC",x"00",x"04",x"05",
															x"02",x"FE",x"FB",x"FB",x"FE",x"03",x"06",x"07",x"04",x"00",x"FD",x"FD",x"00",x"04",x"07",x"06",x"02",x"FE",x"FB",x"FC",x"FF",x"03",x"05",x"03",x"FF",x"FB",x"F9",x"FA",x"FE",x"02",x"04",x"03",x"00",x"FD",x"FB",x"FD",x"02",x"06",x"08",x"06",x"02",x"FE",x"FC",x"FE",x"02",x"05",x"05",x"02",x"FE",x"FB",x"FA",x"FD",x"00",x"03",x"03",x"00",x"FD",x"FA",x"FB",x"FF",x"03",x"06",x"06",x"02",x"FE",x"FC",x"FC",x"FF",x"04",x"05",x"00",x"FC",x"FA",x"F8",x"F7",x"F6",x"FA",x"04",x"10",x"19",x"1E",x"1C",x"14",x"0A",x"FE",x"F4",x"EC",x"E6",x"E1",x"DE",x"DE",x"DF",x"E1",x"E2",x"E5",x"EA",x"F1",x"FA",x"04",x"0E",
															x"15",x"1B",x"1E",x"20",x"21",x"20",x"1C",x"17",x"12",x"0D",x"07",x"00",x"F7",x"EC",x"E1",x"D6",x"CD",x"C6",x"C2",x"C0",x"C0",x"C1",x"C5",x"CB",x"D0",x"D5",x"DB",x"E3",x"ED",x"F9",x"04",x"0E",x"17",x"1D",x"21",x"23",x"24",x"24",x"21",x"1D",x"17",x"11",x"0C",x"05",x"FD",x"F4",x"EB",x"E2",x"DA",x"D4",x"D0",x"CE",x"CE",x"CF",x"D3",x"D8",x"DE",x"E5",x"EC",x"F5",x"FE",x"09",x"15",x"20",x"2A",x"31",x"35",x"36",x"36",x"34",x"30",x"2B",x"25",x"1F",x"19",x"11",x"06",x"FB",x"F0",x"E5",x"DC",x"D6",x"D3",x"D2",x"D3",x"D5",x"D8",x"DD",x"E2",x"E8",x"EE",x"F5",x"FD",x"07",x"12",x"1C",x"24",x"2A",x"2E",x"2F",
															x"30",x"2E",x"2B",x"26",x"20",x"1B",x"14",x"0D",x"04",x"F9",x"ED",x"E2",x"D9",x"D3",x"D0",x"CF",x"D0",x"D2",x"D6",x"DB",x"E1",x"E7",x"EE",x"F6",x"01",x"0C",x"18",x"23",x"2B",x"31",x"35",x"37",x"36",x"34",x"2F",x"29",x"23",x"1D",x"16",x"0D",x"02",x"F6",x"EB",x"E1",x"D9",x"D4",x"D1",x"D0",x"D1",x"D3",x"D8",x"DD",x"E2",x"E8",x"EF",x"F9",x"03",x"0F",x"19",x"23",x"2A",x"2F",x"32",x"32",x"31",x"2D",x"28",x"22",x"1D",x"16",x"0F",x"05",x"FA",x"EF",x"E4",x"DC",x"D5",x"D1",x"CF",x"CF",x"D0",x"D3",x"D8",x"DE",x"E4",x"EB",x"F4",x"FE",x"09",x"14",x"1F",x"28",x"2E",x"32",x"33",x"32",x"2F",x"2B",x"26",x"20",
															x"1B",x"13",x"0A",x"00",x"F5",x"EA",x"E0",x"D8",x"D3",x"D0",x"CE",x"CF",x"D1",x"D6",x"DC",x"E2",x"E9",x"F1",x"FA",x"05",x"10",x"1A",x"24",x"2B",x"2F",x"32",x"32",x"30",x"2C",x"28",x"23",x"1E",x"18",x"10",x"07",x"FC",x"F0",x"E5",x"DD",x"D6",x"D1",x"CF",x"CF",x"D1",x"D5",x"DB",x"E1",x"E7",x"ED",x"F5",x"FE",x"09",x"15",x"1F",x"26",x"2C",x"2F",x"30",x"2F",x"2D",x"29",x"24",x"1F",x"19",x"13",x"0B",x"01",x"F6",x"EB",x"E1",x"D9",x"D3",x"D0",x"CF",x"D0",x"D3",x"D8",x"DE",x"E4",x"EA",x"F1",x"FA",x"04",x"0F",x"1A",x"23",x"2A",x"2F",x"31",x"31",x"30",x"2D",x"29",x"23",x"1D",x"17",x"0F",x"06",x"FB",x"F0",
															x"E5",x"DC",x"D5",x"D1",x"CF",x"CF",x"D1",x"D5",x"DA",x"E0",x"E5",x"EB",x"F3",x"FD",x"08",x"13",x"1D",x"25",x"2C",x"30",x"32",x"32",x"31",x"2D",x"28",x"22",x"1C",x"15",x"0D",x"04",x"F9",x"ED",x"E2",x"DA",x"D4",x"D1",x"CF",x"D0",x"D2",x"D6",x"DB",x"E1",x"E6",x"ED",x"F6",x"00",x"0C",x"17",x"22",x"2A",x"30",x"33",x"34",x"33",x"30",x"2B",x"25",x"1F",x"19",x"12",x"08",x"FD",x"F1",x"E6",x"DC",x"D5",x"D0",x"CE",x"CE",x"CF",x"D3",x"D8",x"DD",x"E3",x"EA",x"F2",x"FC",x"07",x"12",x"1D",x"26",x"2E",x"33",x"35",x"35",x"33",x"2E",x"29",x"23",x"1D",x"17",x"0F",x"05",x"FA",x"EE",x"E3",x"DB",x"D4",x"D0",x"CE",
															x"CD",x"CF",x"D3",x"D9",x"DE",x"E4",x"EB",x"F3",x"FD",x"08",x"14",x"1F",x"27",x"2E",x"31",x"33",x"32",x"30",x"2C",x"27",x"23",x"1D",x"16",x"0E",x"04",x"F9",x"EE",x"E4",x"DC",x"D7",x"D4",x"D2",x"D2",x"D5",x"D9",x"DE",x"E3",x"E9",x"F0",x"F8",x"01",x"0C",x"17",x"21",x"28",x"2D",x"2F",x"30",x"2F",x"2C",x"29",x"24",x"20",x"1A",x"13",x"0A",x"00",x"F5",x"EB",x"E2",x"DB",x"D7",x"D4",x"D4",x"D5",x"D8",x"DC",x"E1",x"E6",x"EC",x"F3",x"FC",x"06",x"11",x"1A",x"22",x"27",x"2A",x"2C",x"2C",x"2B",x"28",x"25",x"21",x"1C",x"16",x"0F",x"06",x"FC",x"F2",x"EA",x"E2",x"DD",x"DA",x"D9",x"D9",x"DB",x"DE",x"E2",x"E6",
															x"EA",x"EF",x"F7",x"00",x"09",x"12",x"1A",x"21",x"25",x"27",x"29",x"29",x"28",x"25",x"21",x"1D",x"18",x"11",x"0A",x"01",x"F8",x"EF",x"E7",x"E1",x"DD",x"DB",x"DA",x"DB",x"DD",x"E0",x"E4",x"E8",x"ED",x"F4",x"FC",x"05",x"0E",x"16",x"1E",x"23",x"27",x"28",x"29",x"28",x"25",x"21",x"1D",x"18",x"13",x"0C",x"05",x"FC",x"F4",x"EC",x"E5",x"E1",x"DE",x"DD",x"DD",x"DE",x"E1",x"E4",x"E8",x"EC",x"F2",x"F8",x"00",x"08",x"10",x"18",x"1E",x"22",x"25",x"26",x"26",x"24",x"20",x"1C",x"18",x"14",x"0F",x"08",x"01",x"F9",x"F1",x"EA",x"E5",x"E2",x"E0",x"DF",x"DF",x"E1",x"E4",x"E7",x"EB",x"F0",x"F5",x"FB",x"03",x"0B",
															x"12",x"18",x"1D",x"20",x"22",x"22",x"21",x"1F",x"1C",x"18",x"15",x"11",x"0C",x"06",x"FF",x"F7",x"F0",x"EB",x"E6",x"E4",x"E2",x"E2",x"E2",x"E5",x"E8",x"EB",x"EF",x"F3",x"F9",x"FF",x"06",x"0D",x"13",x"18",x"1C",x"1E",x"1F",x"1F",x"1D",x"1B",x"19",x"16",x"12",x"0E",x"09",x"03",x"FC",x"F5",x"EF",x"EA",x"E6",x"E4",x"E3",x"E3",x"E4",x"E7",x"EA",x"EE",x"F2",x"F6",x"FB",x"02",x"09",x"0F",x"15",x"19",x"1B",x"1D",x"1D",x"1D",x"1B",x"19",x"16",x"13",x"0F",x"0A",x"05",x"FE",x"F8",x"F1",x"EB",x"E7",x"E4",x"E3",x"E3",x"E4",x"E6",x"E9",x"EC",x"F0",x"F4",x"F9",x"FF",x"06",x"0C",x"12",x"17",x"1A",x"1C",x"1D",
															x"1D",x"1C",x"1A",x"18",x"14",x"11",x"0D",x"07",x"01",x"FA",x"F4",x"EE",x"E9",x"E6",x"E5",x"E4",x"E5",x"E6",x"E9",x"EC",x"EF",x"F3",x"F7",x"FC",x"02",x"09",x"0F",x"14",x"18",x"1B",x"1C",x"1C",x"1C",x"1B",x"18",x"15",x"12",x"0E",x"0A",x"04",x"FE",x"F8",x"F2",x"ED",x"E9",x"E6",x"E5",x"E5",x"E6",x"E8",x"EA",x"ED",x"F0",x"F4",x"F9",x"FE",x"04",x"0A",x"10",x"15",x"19",x"1B",x"1C",x"1D",x"1C",x"1A",x"17",x"14",x"10",x"0C",x"08",x"03",x"FD",x"F7",x"F1",x"ED",x"EA",x"E8",x"E7",x"E7",x"E8",x"EA",x"EC",x"EF",x"F2",x"F5",x"FA",x"FF",x"05",x"0B",x"0F",x"14",x"17",x"18",x"19",x"19",x"18",x"16",x"13",x"11",
															x"0E",x"0A",x"06",x"01",x"FB",x"F6",x"F2",x"EE",x"EC",x"EA",x"EA",x"EA",x"EB",x"ED",x"EF",x"F2",x"F5",x"F8",x"FD",x"02",x"07",x"0C",x"11",x"14",x"16",x"17",x"17",x"16",x"14",x"12",x"0F",x"0D",x"0A",x"07",x"03",x"FE",x"F9",x"F5",x"F1",x"EE",x"ED",x"EC",x"EB",x"EC",x"ED",x"F0",x"F2",x"F4",x"F7",x"FB",x"FF",x"04",x"09",x"0D",x"11",x"13",x"15",x"15",x"15",x"14",x"12",x"10",x"0E",x"0C",x"09",x"05",x"01",x"FC",x"F7",x"F3",x"EF",x"ED",x"EC",x"EB",x"EB",x"EC",x"EE",x"F1",x"F3",x"F6",x"FA",x"FE",x"02",x"07",x"0B",x"0F",x"12",x"13",x"14",x"14",x"14",x"13",x"11",x"0F",x"0D",x"0A",x"06",x"02",x"FE",x"F9",
															x"F4",x"F1",x"EE",x"EC",x"EC",x"EC",x"ED",x"EE",x"F0",x"F3",x"F5",x"F8",x"FC",x"00",x"05",x"0A",x"0D",x"10",x"12",x"13",x"14",x"14",x"13",x"12",x"10",x"0E",x"0B",x"08",x"04",x"00",x"FB",x"F6",x"F3",x"F0",x"EE",x"EE",x"ED",x"EE",x"EF",x"F1",x"F3",x"F6",x"F8",x"FB",x"FE",x"01",x"05",x"09",x"0C",x"0F",x"12",x"13",x"13",x"13",x"13",x"11",x"0F",x"0D",x"0A",x"07",x"03",x"FF",x"FA",x"F5",x"F2",x"F0",x"EE",x"ED",x"EE",x"EF",x"F0",x"F2",x"F4",x"F6",x"F8",x"FA",x"FE",x"02",x"07",x"0B",x"0F",x"11",x"12",x"12",x"12",x"12",x"11",x"0C",x"08",x"08",x"08",x"04",x"FC",x"F5",x"F5",x"F9",x"FC",x"FC",x"F5",x"EB",
															x"E4",x"E4",x"EB",x"F9",x"06",x"0D",x"0A",x"00",x"F2",x"E7",x"E4",x"EA",x"F8",x"09",x"15",x"18",x"11",x"02",x"F3",x"EB",x"ED",x"F7",x"07",x"15",x"19",x"14",x"06",x"F4",x"E5",x"E0",x"E5",x"F2",x"01",x"0B",x"0A",x"FE",x"EB",x"D8",x"CF",x"D0",x"DC",x"ED",x"FC",x"01",x"FA",x"EB",x"DA",x"CE",x"CC",x"D5",x"E4",x"F7",x"04",x"08",x"01",x"F3",x"E3",x"D9",x"DA",x"E5",x"F7",x"09",x"13",x"12",x"08",x"F9",x"ED",x"EA",x"F0",x"FF",x"10",x"1D",x"1F",x"17",x"09",x"F8",x"EE",x"EF",x"F9",x"09",x"18",x"1E",x"19",x"0D",x"FC",x"F0",x"ED",x"F3",x"01",x"10",x"19",x"18",x"0F",x"FF",x"F0",x"E9",x"EC",x"F8",x"07",x"15",
															x"19",x"12",x"04",x"F6",x"EC",x"EB",x"F3",x"00",x"0E",x"17",x"17",x"0F",x"00",x"F0",x"E8",x"E9",x"F3",x"02",x"0F",x"15",x"11",x"05",x"F6",x"EB",x"E9",x"F0",x"FE",x"0E",x"16",x"15",x"0C",x"FD",x"EF",x"EA",x"EE",x"F9",x"08",x"14",x"16",x"0F",x"02",x"F3",x"EB",x"EC",x"F5",x"04",x"11",x"17",x"13",x"07",x"F8",x"ED",x"EB",x"F2",x"FF",x"0E",x"16",x"15",x"0C",x"FE",x"F2",x"ED",x"F1",x"FC",x"0B",x"16",x"18",x"12",x"05",x"F6",x"ED",x"ED",x"F5",x"03",x"10",x"16",x"13",x"09",x"FB",x"F0",x"ED",x"F2",x"FF",x"0D",x"16",x"15",x"0D",x"FE",x"F0",x"EA",x"ED",x"F8",x"07",x"13",x"16",x"10",x"03",x"F4",x"EB",x"EB",
															x"F4",x"02",x"0F",x"14",x"11",x"06",x"F7",x"EC",x"EA",x"F1",x"FE",x"0C",x"15",x"14",x"0B",x"FC",x"F0",x"EB",x"EE",x"F9",x"09",x"14",x"17",x"11",x"04",x"F5",x"EC",x"EC",x"F4",x"02",x"0F",x"16",x"13",x"09",x"FA",x"EF",x"ED",x"F2",x"FF",x"0E",x"17",x"17",x"0E",x"FF",x"F2",x"EC",x"EF",x"F9",x"08",x"14",x"16",x"11",x"04",x"F6",x"EE",x"EE",x"F5",x"03",x"10",x"16",x"12",x"08",x"F9",x"EE",x"EB",x"F1",x"FE",x"0D",x"15",x"15",x"0C",x"FE",x"F1",x"EC",x"EF",x"F9",x"08",x"13",x"16",x"11",x"05",x"F6",x"ED",x"EC",x"F3",x"00",x"0E",x"14",x"13",x"09",x"FB",x"EF",x"EC",x"F1",x"FD",x"0C",x"15",x"15",x"0D",x"FF",
															x"F2",x"EC",x"EE",x"F8",x"06",x"12",x"15",x"0F",x"03",x"F5",x"ED",x"EC",x"F4",x"02",x"0F",x"14",x"11",x"07",x"F9",x"EE",x"EB",x"F1",x"FE",x"0C",x"14",x"14",x"0C",x"FE",x"F2",x"ED",x"F0",x"FA",x"08",x"13",x"16",x"11",x"05",x"F6",x"ED",x"EC",x"F4",x"01",x"0F",x"15",x"13",x"0A",x"FC",x"F0",x"ED",x"F2",x"FE",x"0C",x"15",x"15",x"0E",x"00",x"F3",x"EC",x"EE",x"F8",x"06",x"11",x"14",x"0F",x"04",x"F6",x"ED",x"EC",x"F4",x"01",x"0F",x"15",x"12",x"07",x"F9",x"ED",x"EA",x"F0",x"FD",x"0B",x"14",x"15",x"0C",x"FE",x"F1",x"EC",x"EF",x"F9",x"06",x"12",x"16",x"11",x"05",x"F7",x"ED",x"EB",x"F2",x"FF",x"0E",x"16",
															x"15",x"0C",x"FD",x"F0",x"EC",x"F0",x"FB",x"0A",x"15",x"17",x"11",x"03",x"F4",x"EC",x"ED",x"F6",x"04",x"11",x"16",x"13",x"07",x"F9",x"EE",x"EC",x"F2",x"FF",x"0E",x"16",x"15",x"0C",x"FD",x"F0",x"EB",x"EF",x"FA",x"09",x"14",x"16",x"10",x"03",x"F5",x"EE",x"EF",x"F8",x"05",x"12",x"17",x"14",x"09",x"FB",x"EF",x"EC",x"F2",x"FF",x"0D",x"15",x"15",x"0D",x"00",x"F4",x"EF",x"F2",x"FC",x"0A",x"14",x"17",x"11",x"05",x"F7",x"EF",x"EF",x"F7",x"04",x"10",x"16",x"13",x"08",x"FB",x"F1",x"EE",x"F4",x"FF",x"0C",x"14",x"13",x"0B",x"FE",x"F2",x"ED",x"F1",x"FB",x"09",x"13",x"15",x"10",x"04",x"F7",x"EF",x"F0",x"F8",
															x"04",x"10",x"15",x"13",x"09",x"FC",x"F1",x"EE",x"F3",x"FE",x"0B",x"13",x"14",x"0D",x"01",x"F5",x"F0",x"F2",x"FB",x"08",x"13",x"16",x"11",x"06",x"F9",x"F0",x"F0",x"F7",x"03",x"0E",x"14",x"12",x"09",x"FD",x"F3",x"EF",x"F4",x"FF",x"0B",x"13",x"13",x"0C",x"00",x"F4",x"EE",x"F1",x"FA",x"07",x"11",x"14",x"0F",x"04",x"F7",x"F0",x"F0",x"F7",x"03",x"0E",x"13",x"11",x"08",x"FC",x"F2",x"EE",x"F3",x"FD",x"0A",x"12",x"13",x"0C",x"01",x"F5",x"EF",x"F1",x"FA",x"07",x"11",x"14",x"0F",x"05",x"F8",x"F0",x"F0",x"F6",x"02",x"0D",x"12",x"10",x"08",x"FC",x"F3",x"F0",x"F5",x"FF",x"0A",x"11",x"12",x"0B",x"00",x"F5",
															x"F0",x"F2",x"FA",x"06",x"0F",x"12",x"0E",x"04",x"F9",x"F2",x"F2",x"F8",x"02",x"0C",x"11",x"0F",x"07",x"FC",x"F4",x"F1",x"F5",x"FE",x"09",x"10",x"11",x"0B",x"01",x"F7",x"F1",x"F3",x"FA",x"05",x"0E",x"11",x"0E",x"05",x"FA",x"F3",x"F2",x"F7",x"01",x"0B",x"10",x"0F",x"08",x"FD",x"F4",x"F2",x"F5",x"FE",x"09",x"10",x"10",x"0B",x"01",x"F7",x"F2",x"F3",x"FA",x"05",x"0E",x"10",x"0D",x"04",x"FA",x"F3",x"F3",x"F8",x"01",x"0B",x"0F",x"0E",x"07",x"FD",x"F5",x"F1",x"F5",x"FD",x"07",x"0E",x"10",x"0B",x"01",x"F8",x"F3",x"F4",x"FA",x"04",x"0D",x"10",x"0D",x"05",x"FB",x"F4",x"F3",x"F8",x"00",x"0A",x"0E",x"0D",
															x"07",x"FE",x"F6",x"F3",x"F6",x"FD",x"07",x"0D",x"0E",x"0A",x"01",x"F8",x"F4",x"F5",x"FB",x"04",x"0C",x"0E",x"0C",x"04",x"FB",x"F5",x"F4",x"F8",x"01",x"09",x"0E",x"0D",x"07",x"FE",x"F6",x"F3",x"F6",x"FC",x"05",x"0C",x"0E",x"0A",x"02",x"FA",x"F4",x"F4",x"FA",x"02",x"0A",x"0D",x"0C",x"05",x"FC",x"F6",x"F4",x"F7",x"FF",x"08",x"0D",x"0C",x"07",x"FF",x"F8",x"F4",x"F6",x"FD",x"05",x"0C",x"0D",x"0A",x"02",x"FA",x"F5",x"F6",x"FA",x"02",x"0A",x"0D",x"0B",x"05",x"FC",x"F6",x"F5",x"F9",x"00",x"08",x"0C",x"0B",x"06",x"FF",x"F8",x"F5",x"F7",x"FD",x"04",x"0A",x"0C",x"09",x"02",x"FA",x"F6",x"F6",x"FB",x"02",
															x"09",x"0C",x"0A",x"04",x"FD",x"F7",x"F6",x"F9",x"FF",x"06",x"0A",x"0A",x"06",x"FF",x"F9",x"F6",x"F8",x"FE",x"05",x"0A",x"0B",x"08",x"01",x"FA",x"F7",x"F7",x"FC",x"02",x"09",x"0B",x"09",x"04",x"FD",x"F8",x"F7",x"FA",x"00",x"07",x"0A",x"09",x"05",x"FE",x"F9",x"F6",x"F8",x"FD",x"04",x"09",x"0A",x"08",x"02",x"FB",x"F7",x"F8",x"FC",x"02",x"08",x"0A",x"08",x"03",x"FD",x"F8",x"F7",x"FA",x"00",x"06",x"09",x"09",x"05",x"FF",x"F9",x"F7",x"F9",x"FE",x"05",x"09",x"0A",x"07",x"02",x"FB",x"F7",x"F8",x"FC",x"02",x"08",x"0A",x"08",x"04",x"FD",x"F8",x"F7",x"FA",x"FF",x"05",x"09",x"09",x"05",x"FF",x"F9",x"F7",
															x"F8",x"FD",x"03",x"08",x"0A",x"08",x"02",x"FC",x"F8",x"F8",x"FC",x"02",x"08",x"0A",x"08",x"03",x"FC",x"F7",x"F6",x"F9",x"FE",x"05",x"08",x"08",x"05",x"FF",x"F9",x"F7",x"F8",x"FD",x"04",x"09",x"0A",x"07",x"02",x"FB",x"F7",x"F8",x"FC",x"02",x"08",x"0A",x"08",x"03",x"FD",x"F8",x"F7",x"F9",x"FF",x"05",x"09",x"08",x"05",x"FF",x"FA",x"F7",x"F9",x"FD",x"03",x"08",x"09",x"07",x"02",x"FC",x"F9",x"F9",x"FC",x"01",x"06",x"08",x"07",x"03",x"FD",x"F8",x"F7",x"F9",x"FE",x"03",x"07",x"06",x"04",x"FE",x"FA",x"F8",x"FA",x"FE",x"04",x"08",x"0A",x"07",x"02",x"FC",x"F8",x"F8",x"FB",x"00",x"06",x"09",x"08",x"04",
															x"FF",x"FA",x"F8",x"FA",x"FE",x"03",x"05",x"04",x"01",x"FC",x"F7",x"F3",x"F3",x"F3",x"F7",x"FF",x"0B",x"15",x"1D",x"20",x"1A",x"0C",x"FB",x"EB",x"E0",x"DC",x"E2",x"EC",x"F8",x"02",x"05",x"00",x"F5",x"EA",x"E1",x"DE",x"E2",x"EC",x"F7",x"01",x"06",x"04",x"FB",x"F0",x"E5",x"DF",x"E0",x"EA",x"F9",x"05",x"0E",x"10",x"0A",x"FD",x"EF",x"E2",x"DB",x"DC",x"E4",x"F0",x"FA",x"00",x"FC",x"EE",x"DC",x"CB",x"BD",x"B4",x"B3",x"B9",x"C2",x"CA",x"CF",x"CC",x"C3",x"B6",x"AC",x"A6",x"A8",x"B3",x"C3",x"D4",x"E3",x"EC",x"EE",x"E9",x"E3",x"E0",x"E2",x"EE",x"03",x"1B",x"31",x"43",x"4A",x"48",x"3E",x"32",x"27",x"24",
															x"2B",x"3A",x"49",x"56",x"5B",x"54",x"43",x"2C",x"15",x"03",x"FA",x"FA",x"00",x"07",x"0B",x"07",x"F9",x"E4",x"D1",x"C2",x"BA",x"BD",x"C7",x"D5",x"E2",x"EC",x"EE",x"E8",x"DE",x"D4",x"CF",x"D3",x"E1",x"F7",x"0F",x"25",x"33",x"35",x"2E",x"23",x"17",x"10",x"13",x"1E",x"2F",x"3F",x"4A",x"4A",x"3E",x"2A",x"13",x"FF",x"F3",x"F1",x"F7",x"FF",x"06",x"06",x"FB",x"E9",x"D5",x"C3",x"B9",x"BA",x"C4",x"D2",x"E1",x"EC",x"EE",x"E8",x"DE",x"D5",x"D1",x"D6",x"E7",x"FF",x"18",x"2C",x"38",x"3A",x"33",x"28",x"1E",x"18",x"1D",x"2A",x"3B",x"4B",x"55",x"54",x"47",x"34",x"1D",x"0A",x"FE",x"FD",x"02",x"09",x"0F",x"0D",
															x"00",x"EC",x"D7",x"C5",x"BA",x"BA",x"C3",x"D1",x"DE",x"E7",x"E7",x"E0",x"D5",x"CB",x"C7",x"CD",x"DD",x"F4",x"0D",x"21",x"2E",x"30",x"29",x"1F",x"16",x"12",x"17",x"25",x"37",x"47",x"51",x"4F",x"41",x"2E",x"19",x"08",x"FE",x"FD",x"01",x"08",x"0B",x"09",x"FC",x"E7",x"D2",x"C1",x"B8",x"BA",x"C4",x"D2",x"DE",x"E6",x"E6",x"DE",x"D3",x"CA",x"C8",x"D0",x"E3",x"FB",x"14",x"29",x"35",x"36",x"2F",x"25",x"1D",x"1A",x"21",x"30",x"40",x"4F",x"56",x"53",x"45",x"31",x"1D",x"0C",x"04",x"04",x"09",x"0D",x"0E",x"07",x"F8",x"E3",x"CD",x"BD",x"B6",x"BA",x"C6",x"D3",x"DF",x"E4",x"E2",x"D9",x"CE",x"C7",x"C5",x"CD",
															x"E0",x"F8",x"10",x"24",x"2E",x"2E",x"28",x"20",x"19",x"18",x"1F",x"2D",x"3C",x"4A",x"50",x"4D",x"3F",x"2D",x"1A",x"0C",x"05",x"06",x"0A",x"0E",x"0F",x"08",x"F8",x"E3",x"CF",x"BF",x"B9",x"BE",x"C9",x"D6",x"E1",x"E6",x"E2",x"D7",x"CB",x"C3",x"C3",x"CD",x"E1",x"F8",x"0F",x"21",x"2A",x"29",x"22",x"1B",x"16",x"17",x"20",x"2E",x"3F",x"4C",x"53",x"4F",x"42",x"31",x"1F",x"11",x"0C",x"0D",x"12",x"16",x"16",x"0E",x"FE",x"E9",x"D4",x"C4",x"BE",x"C2",x"CD",x"D9",x"E2",x"E5",x"DF",x"D4",x"C7",x"BE",x"BD",x"C8",x"DC",x"F4",x"0C",x"1E",x"27",x"25",x"1D",x"15",x"10",x"13",x"1E",x"2F",x"41",x"4F",x"55",x"51",
															x"41",x"2D",x"1C",x"0F",x"0A",x"0D",x"13",x"18",x"18",x"0F",x"FE",x"E8",x"D1",x"C0",x"B9",x"BD",x"C9",x"D8",x"E4",x"E8",x"E3",x"D7",x"CA",x"C0",x"BE",x"C7",x"DB",x"F4",x"0D",x"21",x"2A",x"29",x"21",x"18",x"12",x"12",x"1C",x"2B",x"3C",x"4A",x"51",x"4D",x"3F",x"2E",x"1C",x"0F",x"0A",x"0E",x"14",x"19",x"1A",x"12",x"01",x"EB",x"D6",x"C5",x"BE",x"C3",x"D0",x"DC",x"E6",x"E9",x"E4",x"D8",x"CB",x"C2",x"C1",x"CA",x"DD",x"F4",x"0A",x"1D",x"26",x"25",x"1F",x"18",x"13",x"15",x"20",x"2F",x"40",x"4D",x"54",x"50",x"43",x"33",x"23",x"16",x"12",x"15",x"1B",x"1F",x"1E",x"15",x"04",x"EE",x"D8",x"C8",x"C1",x"C5",
															x"D0",x"DC",x"E5",x"E8",x"E1",x"D6",x"CA",x"C2",x"C1",x"CB",x"DE",x"F5",x"0B",x"1C",x"24",x"23",x"1D",x"18",x"15",x"18",x"23",x"31",x"40",x"4C",x"51",x"4C",x"40",x"30",x"21",x"15",x"11",x"13",x"17",x"19",x"18",x"0F",x"FF",x"EC",x"D9",x"CB",x"C5",x"C8",x"D2",x"DC",x"E5",x"E7",x"E3",x"D9",x"CF",x"C9",x"C9",x"D2",x"E3",x"F7",x"0A",x"19",x"20",x"1F",x"1A",x"14",x"12",x"15",x"1E",x"2B",x"37",x"41",x"44",x"3F",x"34",x"27",x"1A",x"12",x"10",x"12",x"16",x"19",x"17",x"0E",x"00",x"F0",x"E0",x"D4",x"CF",x"D3",x"DC",x"E6",x"EE",x"F0",x"EB",x"E1",x"D8",x"D1",x"D0",x"D8",x"E6",x"F6",x"07",x"13",x"19",x"18",
															x"14",x"10",x"0E",x"11",x"19",x"24",x"2E",x"37",x"3A",x"37",x"2F",x"25",x"1B",x"14",x"12",x"15",x"18",x"19",x"17",x"0F",x"02",x"F3",x"E5",x"DB",x"D7",x"DA",x"E0",x"E8",x"ED",x"EC",x"E6",x"DD",x"D5",x"D0",x"D1",x"D9",x"E5",x"F4",x"02",x"0D",x"12",x"12",x"0F",x"0D",x"0C",x"10",x"18",x"22",x"2C",x"33",x"36",x"33",x"2B",x"22",x"19",x"13",x"12",x"13",x"16",x"18",x"16",x"0F",x"03",x"F5",x"E8",x"DE",x"DB",x"DD",x"E3",x"EA",x"EF",x"EF",x"EA",x"E2",x"DB",x"D6",x"D6",x"DD",x"EA",x"F8",x"05",x"0E",x"12",x"11",x"0E",x"0B",x"0B",x"0F",x"18",x"21",x"2A",x"30",x"32",x"2E",x"26",x"1D",x"14",x"0F",x"0E",x"11",
															x"14",x"15",x"13",x"0C",x"00",x"F3",x"E7",x"DE",x"DB",x"DF",x"E5",x"ED",x"F2",x"F1",x"EC",x"E3",x"DC",x"D7",x"D8",x"E0",x"EC",x"FA",x"07",x"0F",x"12",x"0F",x"0B",x"08",x"07",x"0D",x"16",x"21",x"2A",x"30",x"30",x"2A",x"22",x"19",x"11",x"0E",x"10",x"15",x"19",x"1A",x"17",x"0D",x"00",x"F2",x"E6",x"DF",x"DE",x"E3",x"EB",x"F1",x"F5",x"F3",x"EC",x"E2",x"D9",x"D5",x"D7",x"E0",x"ED",x"FA",x"05",x"0C",x"0C",x"09",x"05",x"02",x"04",x"0B",x"16",x"21",x"29",x"2E",x"2D",x"27",x"1E",x"16",x"11",x"0F",x"13",x"17",x"1B",x"1B",x"17",x"0D",x"00",x"F3",x"E8",x"E1",x"E1",x"E6",x"ED",x"F3",x"F6",x"F3",x"EC",x"E3",
															x"DB",x"D8",x"DB",x"E3",x"EF",x"FC",x"06",x"0C",x"0D",x"0B",x"08",x"05",x"06",x"0B",x"14",x"1C",x"24",x"29",x"28",x"24",x"1C",x"14",x"0E",x"0B",x"0D",x"10",x"14",x"15",x"12",x"0A",x"FF",x"F4",x"EB",x"E5",x"E4",x"E8",x"ED",x"F2",x"F5",x"F3",x"ED",x"E6",x"E0",x"DD",x"DF",x"E6",x"F0",x"FA",x"03",x"08",x"09",x"07",x"04",x"02",x"03",x"09",x"12",x"1B",x"22",x"26",x"25",x"20",x"19",x"13",x"0E",x"0D",x"0F",x"13",x"15",x"16",x"13",x"0B",x"01",x"F6",x"EE",x"E9",x"E9",x"ED",x"F2",x"F6",x"F8",x"F5",x"EF",x"E8",x"E1",x"DE",x"E1",x"E8",x"F1",x"FA",x"02",x"05",x"05",x"03",x"00",x"00",x"02",x"09",x"11",x"1A",
															x"20",x"22",x"20",x"1C",x"16",x"11",x"0E",x"0E",x"10",x"14",x"17",x"16",x"12",x"0A",x"00",x"F6",x"EF",x"EA",x"EA",x"EE",x"F3",x"F6",x"F8",x"F5",x"EF",x"E8",x"E2",x"DF",x"E1",x"E7",x"F0",x"FA",x"01",x"05",x"05",x"03",x"00",x"FF",x"01",x"07",x"0E",x"16",x"1C",x"1F",x"1D",x"18",x"13",x"0E",x"0B",x"0C",x"0E",x"11",x"13",x"13",x"0F",x"08",x"FF",x"F6",x"F0",x"ED",x"EE",x"F1",x"F5",x"F9",x"FA",x"F6",x"F0",x"EA",x"E6",x"E3",x"E6",x"EC",x"F3",x"FA",x"00",x"03",x"03",x"01",x"FF",x"FE",x"01",x"07",x"0E",x"14",x"19",x"1C",x"1A",x"17",x"12",x"0E",x"0B",x"0B",x"0D",x"10",x"12",x"13",x"10",x"0A",x"02",x"FA",
															x"F2",x"EE",x"EE",x"F0",x"F4",x"F7",x"F8",x"F6",x"F1",x"EC",x"E7",x"E5",x"E7",x"EC",x"F3",x"FA",x"FF",x"01",x"00",x"FE",x"FD",x"FD",x"FD",x"03",x"0E",x"16",x"18",x"16",x"15",x"15",x"16",x"14",x"0F",x"0A",x"09",x"0B",x"11",x"18",x"1A",x"14",x"06",x"F2",x"E0",x"D5",x"D5",x"DE",x"EC",x"FA",x"00",x"FC",x"F1",x"E3",x"D9",x"D9",x"E3",x"F3",x"04",x"10",x"12",x"0C",x"00",x"F5",x"EF",x"F3",x"FE",x"0E",x"1A",x"1E",x"18",x"0B",x"FB",x"F0",x"EE",x"F3",x"FE",x"0A",x"11",x"0E",x"03",x"F4",x"E5",x"DE",x"E1",x"EA",x"F7",x"04",x"09",x"05",x"F9",x"EA",x"DC",x"D8",x"DD",x"EA",x"FB",x"08",x"0C",x"06",x"F9",x"EA",
															x"E2",x"E4",x"EE",x"FF",x"0E",x"16",x"14",x"0A",x"FB",x"EF",x"EC",x"F2",x"FF",x"0E",x"18",x"19",x"11",x"02",x"F4",x"EC",x"EE",x"F8",x"07",x"13",x"18",x"13",x"06",x"F7",x"EC",x"EA",x"F1",x"FF",x"0D",x"15",x"14",x"0A",x"FC",x"F0",x"EB",x"F0",x"FC",x"0B",x"17",x"1A",x"14",x"08",x"F8",x"EC",x"E9",x"F0",x"FD",x"0D",x"16",x"16",x"0D",x"FF",x"F1",x"EB",x"EF",x"FA",x"09",x"15",x"18",x"11",x"03",x"F4",x"EB",x"EC",x"F5",x"03",x"10",x"15",x"11",x"05",x"F6",x"EB",x"E9",x"F0",x"FD",x"0C",x"14",x"13",x"0A",x"FB",x"EE",x"E9",x"EE",x"F9",x"08",x"13",x"15",x"0F",x"03",x"F5",x"ED",x"EF",x"F8",x"06",x"13",x"18",
															x"15",x"0A",x"FB",x"EF",x"EC",x"F1",x"FD",x"0C",x"15",x"15",x"0D",x"00",x"F2",x"EC",x"EE",x"F9",x"08",x"14",x"17",x"12",x"05",x"F6",x"EC",x"EB",x"F3",x"01",x"0F",x"15",x"13",x"08",x"F9",x"ED",x"EA",x"EF",x"FC",x"0B",x"14",x"14",x"0C",x"FD",x"EF",x"E8",x"EB",x"F6",x"05",x"12",x"15",x"0F",x"03",x"F4",x"EB",x"EB",x"F3",x"01",x"0F",x"16",x"14",x"09",x"FA",x"ED",x"E9",x"EE",x"FA",x"09",x"14",x"15",x"0E",x"00",x"F2",x"EB",x"ED",x"F7",x"07",x"13",x"17",x"12",x"06",x"F7",x"ED",x"EC",x"F3",x"01",x"10",x"17",x"15",x"0A",x"FB",x"EE",x"EA",x"F0",x"FC",x"0B",x"15",x"15",x"0D",x"FF",x"F1",x"EA",x"ED",x"F7",
															x"06",x"12",x"16",x"11",x"04",x"F5",x"EB",x"EB",x"F3",x"01",x"10",x"17",x"14",x"0A",x"FB",x"EE",x"E9",x"EE",x"FA",x"09",x"14",x"15",x"0E",x"01",x"F2",x"EB",x"EC",x"F6",x"05",x"12",x"17",x"12",x"06",x"F7",x"EC",x"EA",x"F2",x"00",x"0E",x"15",x"14",x"0A",x"FB",x"EE",x"EA",x"EE",x"FA",x"0A",x"14",x"15",x"0E",x"00",x"F1",x"EA",x"EB",x"F5",x"05",x"12",x"16",x"12",x"05",x"F6",x"EC",x"EB",x"F3",x"00",x"0F",x"16",x"15",x"0C",x"FD",x"F0",x"EA",x"EE",x"F9",x"09",x"14",x"16",x"10",x"02",x"F2",x"EA",x"EB",x"F5",x"04",x"12",x"18",x"14",x"08",x"F8",x"ED",x"EA",x"F1",x"FF",x"0D",x"16",x"15",x"0B",x"FC",x"EF",
															x"EA",x"EE",x"FA",x"09",x"14",x"16",x"0F",x"01",x"F2",x"EA",x"EB",x"F5",x"04",x"11",x"16",x"12",x"06",x"F6",x"EC",x"EB",x"F3",x"00",x"0E",x"15",x"13",x"0B",x"FD",x"F0",x"EB",x"EE",x"F8",x"07",x"13",x"16",x"10",x"03",x"F5",x"EC",x"EC",x"F4",x"02",x"10",x"16",x"13",x"09",x"FB",x"EF",x"EC",x"F1",x"FD",x"0B",x"14",x"14",x"0C",x"FE",x"F1",x"EC",x"EF",x"F9",x"08",x"13",x"15",x"10",x"04",x"F6",x"ED",x"EE",x"F6",x"03",x"0F",x"15",x"12",x"08",x"FA",x"F0",x"EE",x"F4",x"00",x"0D",x"14",x"14",x"0D",x"01",x"F5",x"EF",x"F1",x"FA",x"07",x"11",x"15",x"11",x"06",x"F9",x"F0",x"EF",x"F6",x"02",x"0E",x"14",x"12",
															x"0A",x"FD",x"F3",x"F0",x"F4",x"FE",x"0A",x"12",x"12",x"0C",x"00",x"F5",x"EF",x"F1",x"FA",x"07",x"10",x"13",x"0F",x"05",x"F8",x"F1",x"F0",x"F7",x"02",x"0D",x"12",x"10",x"08",x"FC",x"F3",x"F1",x"F5",x"FF",x"0A",x"12",x"13",x"0D",x"02",x"F6",x"F0",x"F1",x"F9",x"05",x"0F",x"13",x"10",x"06",x"FA",x"F1",x"F0",x"F6",x"01",x"0C",x"12",x"11",x"0A",x"FE",x"F4",x"F1",x"F4",x"FE",x"09",x"11",x"12",x"0C",x"01",x"F6",x"F0",x"F2",x"FA",x"06",x"0F",x"12",x"0E",x"05",x"F9",x"F2",x"F1",x"F7",x"01",x"0C",x"11",x"0F",x"07",x"FC",x"F3",x"F1",x"F6",x"FF",x"0A",x"11",x"11",x"0B",x"01",x"F6",x"F1",x"F2",x"FA",x"05",
															x"0E",x"11",x"0E",x"05",x"F9",x"F2",x"F1",x"F7",x"01",x"0C",x"11",x"10",x"08",x"FD",x"F4",x"F1",x"F5",x"FE",x"08",x"10",x"10",x"0A",x"00",x"F6",x"F1",x"F3",x"FA",x"05",x"0E",x"11",x"0D",x"04",x"FA",x"F3",x"F2",x"F8",x"01",x"0B",x"10",x"0E",x"07",x"FD",x"F5",x"F2",x"F6",x"FF",x"09",x"0F",x"10",x"0A",x"01",x"F7",x"F2",x"F3",x"FA",x"04",x"0D",x"10",x"0E",x"06",x"FB",x"F4",x"F2",x"F7",x"00",x"0A",x"0F",x"0F",x"08",x"FF",x"F6",x"F3",x"F5",x"FC",x"06",x"0D",x"0F",x"0A",x"02",x"F8",x"F3",x"F3",x"F9",x"03",x"0C",x"0F",x"0D",x"05",x"FB",x"F4",x"F3",x"F7",x"00",x"09",x"0E",x"0D",x"07",x"FE",x"F6",x"F3",
															x"F6",x"FD",x"07",x"0E",x"0E",x"0A",x"01",x"F8",x"F3",x"F4",x"F9",x"03",x"0B",x"0F",x"0C",x"06",x"FC",x"F5",x"F3",x"F7",x"FF",x"08",x"0D",x"0D",x"08",x"FF",x"F7",x"F4",x"F5",x"FC",x"05",x"0C",x"0E",x"0A",x"02",x"F9",x"F4",x"F4",x"F9",x"02",x"0B",x"0E",x"0C",x"06",x"FD",x"F5",x"F3",x"F7",x"FF",x"08",x"0D",x"0D",x"08",x"FF",x"F7",x"F3",x"F6",x"FC",x"05",x"0C",x"0E",x"0A",x"02",x"F9",x"F3",x"F3",x"F8",x"01",x"0A",x"0E",x"0D",x"07",x"FD",x"F5",x"F3",x"F6",x"FE",x"07",x"0D",x"0D",x"09",x"00",x"F8",x"F4",x"F5",x"FB",x"04",x"0B",x"0E",x"0A",x"03",x"FA",x"F4",x"F3",x"F8",x"01",x"0A",x"0E",x"0C",x"06",
															x"FD",x"F6",x"F4",x"F7",x"FE",x"07",x"0C",x"0C",x"08",x"00",x"F8",x"F4",x"F6",x"FC",x"05",x"0C",x"0D",x"0A",x"02",x"F9",x"F4",x"F4",x"F9",x"01",x"0A",x"0D",x"0C",x"06",x"FD",x"F6",x"F4",x"F7",x"FE",x"06",x"0C",x"0C",x"08",x"00",x"F8",x"F4",x"F6",x"FC",x"04",x"0A",x"0C",x"09",x"02",x"FA",x"F5",x"F5",x"F9",x"01",x"09",x"0C",x"0B",x"05",x"FD",x"F7",x"F5",x"F8",x"FF",x"06",x"0B",x"0B",x"07",x"FF",x"F8",x"F5",x"F7",x"FD",x"04",x"0A",x"0C",x"08",x"02",x"FA",x"F5",x"F5",x"FA",x"01",x"08",x"0C",x"0A",x"05",x"FD",x"F7",x"F5",x"F8",x"FE",x"06",x"0A",x"0B",x"07",x"00",x"F9",x"F6",x"F7",x"FC",x"03",x"09",
															x"0B",x"08",x"02",x"FB",x"F6",x"F6",x"FA",x"01",x"07",x"0B",x"0A",x"05",x"FE",x"F8",x"F6",x"F9",x"FF",x"05",x"0A",x"0A",x"06",x"00",x"F9",x"F6",x"F7",x"FC",x"03",x"09",x"0B",x"08",x"02",x"FB",x"F6",x"F6",x"FA",x"00",x"07",x"0B",x"0A",x"05",x"FE",x"F9",x"F6",x"F9",x"FE",x"05",x"0A",x"0A",x"07",x"00",x"FA",x"F6",x"F7",x"FC",x"03",x"09",x"0B",x"09",x"03",x"FC",x"F7",x"F7",x"FA",x"00",x"06",x"09",x"09",x"05",x"FF",x"F9",x"F7",x"F9",x"FE",x"05",x"09",x"09",x"06",x"00",x"FA",x"F7",x"F7",x"FC",x"02",x"06",x"08",x"06",x"01",x"FC",x"F8",x"F8",x"FB",x"01",x"07",x"0B",x"0B",x"07",x"01",x"FA",x"F7",x"F8",
															x"FC",x"02",x"07",x"08",x"06",x"01",x"FC",x"F8",x"F8",x"FB",x"01",x"06",x"08",x"06",x"02",x"FD",x"F9",x"F8",x"FA",x"FF",x"04",x"06",x"05",x"02",x"FC",x"F8",x"F7",x"FA",x"FF",x"05",x"09",x"09",x"05",x"FF",x"F9",x"F6",x"F7",x"FA",x"00",x"05",x"05",x"01",x"FC",x"F5",x"F0",x"EF",x"F0",x"F3",x"F9",x"01",x"0C",x"16",x"1B",x"1B",x"15",x"09",x"F8",x"E8",x"DC",x"D6",x"D7",x"DF",x"ED",x"FB",x"05",x"09",x"07",x"FE",x"F2",x"E7",x"E1",x"DF",x"E3",x"ED",x"F9",x"02",x"07",x"07",x"01",x"F6",x"E8",x"DC",x"D4",x"D2",x"D6",x"E1",x"EF",x"FB",x"01",x"01",x"FA",x"ED",x"DC",x"CC",x"C1",x"BB",x"BE",x"C8",x"D5",x"E0",
															x"E7",x"E7",x"E2",x"D6",x"C6",x"B8",x"AE",x"A8",x"A8",x"B0",x"BD",x"CA",x"D5",x"DB",x"DC",x"D6",x"CC",x"C5",x"C3",x"C7",x"D1",x"E1",x"F5",x"06",x"14",x"1C",x"1D",x"18",x"11",x"0C",x"0B",x"0F",x"1A",x"2B",x"3E",x"4C",x"56",x"59",x"53",x"47",x"38",x"2A",x"20",x"1B",x"1D",x"25",x"2E",x"34",x"36",x"30",x"23",x"11",x"FC",x"EA",x"DE",x"D8",x"D8",x"DD",x"E4",x"E8",x"EA",x"E7",x"E0",x"D4",x"C7",x"BE",x"BB",x"BE",x"C8",x"D7",x"E7",x"F5",x"FF",x"04",x"02",x"FC",x"F5",x"F2",x"F3",x"FB",x"09",x"1C",x"2F",x"3D",x"45",x"46",x"3E",x"31",x"23",x"17",x"10",x"0F",x"16",x"22",x"2C",x"32",x"32",x"29",x"19",x"04",
															x"F1",x"E2",x"D9",x"D7",x"DC",x"E5",x"EC",x"F0",x"EE",x"E7",x"DA",x"CD",x"C4",x"C1",x"C3",x"CD",x"DD",x"ED",x"FC",x"06",x"0B",x"0B",x"04",x"FE",x"FA",x"FA",x"00",x"0E",x"22",x"35",x"45",x"50",x"52",x"4C",x"3F",x"30",x"23",x"1A",x"16",x"1B",x"26",x"30",x"37",x"37",x"2F",x"1F",x"09",x"F4",x"E2",x"D6",x"D1",x"D5",x"DC",x"E3",x"E7",x"E7",x"DF",x"D1",x"C2",x"B7",x"B1",x"B3",x"BC",x"CB",x"DE",x"EE",x"FA",x"00",x"00",x"FA",x"F3",x"F0",x"F2",x"FA",x"0A",x"1F",x"34",x"46",x"51",x"54",x"4D",x"40",x"31",x"24",x"1C",x"19",x"1E",x"29",x"33",x"39",x"39",x"31",x"20",x"0B",x"F6",x"E5",x"D9",x"D5",x"D9",x"E2",
															x"E8",x"EC",x"EB",x"E5",x"D8",x"C9",x"BE",x"B9",x"BA",x"C3",x"D4",x"E6",x"F5",x"00",x"06",x"05",x"FD",x"F6",x"F2",x"F3",x"FA",x"09",x"1E",x"33",x"42",x"4B",x"4D",x"47",x"3A",x"2B",x"1F",x"16",x"13",x"18",x"22",x"2C",x"33",x"34",x"2E",x"1E",x"09",x"F4",x"E3",x"D7",x"D3",x"D8",x"E0",x"E8",x"EC",x"EC",x"E6",x"D8",x"C9",x"BD",x"B7",x"B9",x"C3",x"D4",x"E6",x"F5",x"00",x"05",x"03",x"FB",x"F3",x"EF",x"F0",x"F7",x"06",x"1C",x"31",x"41",x"4A",x"4C",x"45",x"37",x"29",x"1D",x"16",x"14",x"1A",x"26",x"31",x"38",x"38",x"31",x"21",x"0B",x"F5",x"E5",x"DA",x"D6",x"DB",x"E5",x"ED",x"F1",x"EF",x"E8",x"DA",x"CA",
															x"BD",x"B7",x"B8",x"C2",x"D3",x"E6",x"F7",x"02",x"07",x"04",x"FB",x"F1",x"EC",x"ED",x"F5",x"04",x"1A",x"30",x"41",x"4B",x"4D",x"45",x"37",x"29",x"1D",x"16",x"16",x"1C",x"28",x"33",x"3A",x"38",x"31",x"20",x"09",x"F4",x"E5",x"DC",x"D9",x"DC",x"E4",x"EB",x"ED",x"EB",x"E4",x"D6",x"C6",x"B9",x"B4",x"B6",x"BF",x"D0",x"E3",x"F4",x"FF",x"03",x"01",x"F9",x"F1",x"ED",x"EF",x"F7",x"07",x"1C",x"30",x"40",x"4A",x"4C",x"47",x"3B",x"2F",x"25",x"1F",x"1E",x"22",x"2B",x"33",x"37",x"37",x"30",x"21",x"0D",x"FB",x"ED",x"E4",x"DF",x"E1",x"E7",x"EB",x"ED",x"EA",x"E2",x"D6",x"C9",x"BF",x"BA",x"BC",x"C4",x"D2",x"E2",
															x"F0",x"FA",x"00",x"00",x"FC",x"F7",x"F5",x"F6",x"FD",x"09",x"1B",x"2C",x"3B",x"45",x"49",x"46",x"3E",x"34",x"2B",x"24",x"21",x"23",x"28",x"2E",x"33",x"33",x"2E",x"22",x"13",x"03",x"F5",x"EA",x"E4",x"E4",x"E8",x"EB",x"ED",x"EB",x"E6",x"DD",x"D1",x"C8",x"C3",x"C3",x"CA",x"D6",x"E5",x"F1",x"FA",x"00",x"00",x"FC",x"F8",x"F5",x"F7",x"FC",x"07",x"16",x"26",x"34",x"3E",x"43",x"41",x"39",x"30",x"27",x"21",x"1D",x"1E",x"24",x"29",x"2D",x"2E",x"2A",x"20",x"12",x"03",x"F6",x"EC",x"E7",x"E8",x"EB",x"EF",x"F0",x"EE",x"E9",x"DF",x"D4",x"CB",x"C6",x"C6",x"CC",x"D7",x"E5",x"F0",x"F9",x"FD",x"FD",x"F9",x"F4",
															x"F2",x"F3",x"F9",x"03",x"11",x"21",x"2D",x"36",x"3A",x"38",x"31",x"29",x"23",x"1E",x"1C",x"1E",x"23",x"28",x"2C",x"2D",x"29",x"20",x"14",x"06",x"FB",x"F2",x"ED",x"EC",x"EF",x"F2",x"F3",x"F2",x"ED",x"E4",x"DA",x"D0",x"CA",x"C9",x"CE",x"D7",x"E3",x"EE",x"F6",x"FB",x"FB",x"F7",x"F3",x"F0",x"F1",x"F6",x"00",x"0E",x"1C",x"27",x"2F",x"33",x"32",x"2C",x"25",x"1F",x"1C",x"1B",x"1D",x"22",x"27",x"2A",x"2A",x"26",x"1D",x"11",x"05",x"FA",x"F2",x"EE",x"EE",x"F0",x"F3",x"F4",x"F3",x"EF",x"E7",x"DE",x"D6",x"D1",x"D0",x"D4",x"DD",x"E9",x"F3",x"FA",x"FE",x"FF",x"FB",x"F7",x"F4",x"F4",x"F7",x"FF",x"0B",x"17",
															x"22",x"29",x"2C",x"2B",x"25",x"1F",x"19",x"16",x"14",x"16",x"1A",x"1F",x"22",x"22",x"1F",x"17",x"0D",x"02",x"FA",x"F4",x"F1",x"F2",x"F5",x"F8",x"F9",x"F8",x"F3",x"ED",x"E4",x"DD",x"D8",x"D7",x"DA",x"E2",x"EC",x"F5",x"FC",x"FF",x"FF",x"FB",x"F7",x"F4",x"F4",x"F7",x"FD",x"08",x"13",x"1C",x"23",x"26",x"25",x"20",x"1A",x"15",x"12",x"11",x"13",x"17",x"1B",x"1E",x"1F",x"1D",x"17",x"0E",x"05",x"FD",x"F8",x"F5",x"F5",x"F8",x"FA",x"FB",x"FA",x"F5",x"EE",x"E6",x"DF",x"DB",x"DA",x"DD",x"E4",x"ED",x"F5",x"FA",x"FD",x"FC",x"F9",x"F4",x"F0",x"F0",x"F3",x"F9",x"03",x"0E",x"17",x"1E",x"21",x"21",x"1D",x"18",
															x"14",x"11",x"11",x"13",x"17",x"1C",x"1F",x"20",x"1F",x"19",x"11",x"08",x"01",x"FB",x"F8",x"F8",x"FA",x"FC",x"FD",x"FC",x"F8",x"F1",x"E8",x"E1",x"DC",x"DA",x"DC",x"E2",x"EB",x"F3",x"F8",x"FB",x"FB",x"F7",x"F2",x"EF",x"EF",x"F2",x"F8",x"02",x"0C",x"16",x"1C",x"20",x"21",x"1D",x"19",x"14",x"12",x"11",x"12",x"16",x"1B",x"1E",x"1F",x"1D",x"18",x"10",x"07",x"00",x"FA",x"F7",x"F6",x"F8",x"FB",x"FB",x"FA",x"F7",x"F1",x"E9",x"E3",x"DE",x"DC",x"DE",x"E4",x"EC",x"F3",x"F9",x"FC",x"FC",x"F9",x"F6",x"F3",x"F3",x"F5",x"FB",x"04",x"0D",x"16",x"1B",x"1E",x"1F",x"1C",x"17",x"14",x"11",x"11",x"12",x"15",x"19",
															x"1B",x"1C",x"1A",x"15",x"0D",x"05",x"FE",x"F9",x"F6",x"F6",x"F9",x"FB",x"FC",x"FB",x"F7",x"F1",x"EA",x"E4",x"E0",x"DF",x"E0",x"E6",x"ED",x"F4",x"FA",x"FD",x"FD",x"FA",x"F7",x"F4",x"F4",x"F6",x"FB",x"03",x"0C",x"13",x"19",x"1C",x"1C",x"19",x"15",x"11",x"0F",x"0E",x"10",x"13",x"16",x"18",x"18",x"17",x"12",x"0C",x"05",x"FF",x"FB",x"F8",x"F7",x"F9",x"FB",x"FC",x"FB",x"F9",x"F4",x"ED",x"E8",x"E4",x"E2",x"E3",x"E8",x"EE",x"F5",x"F9",x"FC",x"FC",x"FA",x"F6",x"F5",x"F5",x"F7",x"FC",x"02",x"0A",x"11",x"16",x"19",x"19",x"16",x"13",x"0F",x"0E",x"0E",x"0F",x"12",x"15",x"16",x"16",x"15",x"11",x"0B",x"05",
															x"00",x"FC",x"F9",x"F9",x"FB",x"FD",x"FD",x"FC",x"F9",x"F4",x"EE",x"E9",x"E5",x"E4",x"E4",x"E8",x"EE",x"F5",x"F9",x"FD",x"FD",x"FB",x"F8",x"F6",x"F5",x"F6",x"FA",x"00",x"07",x"0E",x"13",x"15",x"16",x"13",x"10",x"0D",x"0C",x"0D",x"0F",x"13",x"17",x"19",x"1A",x"18",x"14",x"0E",x"07",x"01",x"FD",x"FA",x"FA",x"FB",x"FD",x"FD",x"FD",x"F9",x"F0",x"E9",x"E5",x"E1",x"DA",x"D7",x"D9",x"E4",x"F3",x"02",x"0C",x"11",x"11",x"0D",x"06",x"00",x"FA",x"F5",x"F2",x"EF",x"EE",x"EC",x"EA",x"E8",x"E7",x"E8",x"EA",x"ED",x"F1",x"F4",x"F8",x"FC",x"00",x"04",x"07",x"09",x"0A",x"0B",x"0B",x"0B",x"08",x"04",x"00",x"FC",
															x"F8",x"F3",x"ED",x"E6",x"DF",x"D7",x"CF",x"C7",x"BE",x"B5",x"AD",x"A6",x"A0",x"9B",x"98",x"96",x"96",x"99",x"9D",x"A0",x"A3",x"A6",x"A9",x"AD",x"B3",x"BA",x"C4",x"CE",x"D9",x"E5",x"F1",x"FD",x"08",x"13",x"1E",x"28",x"30",x"35",x"3A",x"3D",x"3F",x"42",x"43",x"44",x"45",x"44",x"41",x"3C",x"36",x"2F",x"27",x"1E",x"14",x"0B",x"02",x"F9",x"F1",x"EA",x"E5",x"E2",x"DF",x"DD",x"DB",x"D8",x"D5",x"D3",x"D3",x"D4",x"D8",x"DD",x"E3",x"EA",x"F2",x"FA",x"03",x"0C",x"14",x"1C",x"23",x"28",x"2B",x"2D",x"2E",x"2E",x"2E",x"2F",x"30",x"2F",x"2C",x"29",x"23",x"1C",x"14",x"0B",x"03",x"FA",x"F1",x"E9",x"E2",x"DB");

	constant Wrecking_Crew_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"03", x"07", x"0F", x"0F", x"3F", x"0E", x"3B", x"00", x"03", x"07", x"0F", x"0F", x"3F", x"01", x"04", x"00", x"80", x"C0", x"E0", x"E0", x"F0", x"00", x"60", x"00", x"80", x"C0", x"A0", x"E0", x"F0", x"E0", x"90", x"77", x"02", x"1F", x"0F", x"07", x"0D", x"1F", x"7F", x"08", x"3D", x"00", x"00", x"05", x"02", x"14", x"14", x"60", x"C0", x"C0", x"CE", x"E0", x"00", x"F0", x"FE", x"90", x"30", x"2E", x"0E", x"8E", x"FF", x"4E", x"4E", x"7F", x"7B", x"1F", x"0F", x"01", x"01", x"00", x"00", x"1E", x"1F", x"1F", x"0F", x"0F", x"1F", x"01", x"03", x"F0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"CE", x"80", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"00", x"03", x"07", x"0F", x"0F", x"00", x"0F", x"3F", x"00", x"03", x"07", x"0F", x"0F", x"3F", x"0F", x"0E", x"00", x"80", x"C0", x"E0", x"E0", x"00", x"C0", x"60", x"00", x"80", x"C0", x"A0", x"E0", x"E0", x"B0", x"80", 
															x"77", x"02", x"1F", x"0F", x"67", x"6D", x"7F", x"7F", x"08", x"3D", x"00", x"00", x"05", x"02", x"14", x"74", x"7F", x"0A", x"00", x"00", x"07", x"0D", x"1F", x"7F", x"00", x"15", x"1F", x"0F", x"05", x"02", x"14", x"14", x"3F", x"1B", x"1F", x"0F", x"0F", x"00", x"00", x"00", x"06", x"1F", x"1F", x"0F", x"0F", x"07", x"0F", x"00", x"F0", x"E0", x"F0", x"F8", x"78", x"00", x"00", x"00", x"CE", x"80", x"FC", x"FE", x"7A", x"00", x"00", x"00", x"40", x"00", x"00", x"4E", x"E0", x"00", x"F0", x"FE", x"B0", x"E0", x"CE", x"8E", x"8E", x"FF", x"4E", x"4E", x"67", x"6A", x"1F", x"0F", x"01", x"01", x"00", x"00", x"1E", x"1F", x"1F", x"0F", x"0F", x"1F", x"01", x"03", x"EE", x"05", x"3F", x"5F", x"EF", x"FD", x"FF", x"7F", x"11", x"7A", x"00", x"00", x"0B", x"12", x"34", x"64", x"C0", x"80", x"80", x"8E", x"E0", x"00", x"F0", x"FE", x"20", x"60", x"4E", x"0E", x"0E", x"FF", x"4E", x"4E", 
															x"1F", x"1B", x"3F", x"3F", x"1F", x"01", x"00", x"00", x"06", x"1F", x"BF", x"FF", x"7F", x"21", x"00", x"00", x"F0", x"E0", x"E0", x"E0", x"F0", x"E0", x"00", x"00", x"CE", x"80", x"E0", x"E0", x"F8", x"F8", x"18", x"30", x"03", x"1F", x"3F", x"3F", x"3F", x"30", x"30", x"30", x"03", x"07", x"0F", x"3F", x"1F", x"0F", x"0F", x"0F", x"80", x"C0", x"E0", x"E0", x"F0", x"10", x"10", x"10", x"80", x"C0", x"A0", x"E0", x"F0", x"E0", x"E0", x"E0", x"38", x"3C", x"1F", x"0F", x"0F", x"1F", x"1F", x"1F", x"0F", x"0B", x"08", x"08", x"0C", x"1F", x"1F", x"1F", x"20", x"7E", x"E0", x"E4", x"E0", x"FE", x"E0", x"F0", x"FE", x"BE", x"3E", x"3E", x"7E", x"FE", x"FE", x"F0", x"1C", x"1C", x"1E", x"1E", x"08", x"08", x"08", x"00", x"1C", x"1C", x"1E", x"1E", x"0E", x"0F", x"0F", x"0F", x"70", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"70", x"F0", x"E0", x"F0", x"00", x"00", x"00", x"00", 
															x"03", x"07", x"0F", x"0F", x"1F", x"10", x"10", x"10", x"03", x"07", x"0F", x"0F", x"1F", x"0F", x"0F", x"0F", x"F0", x"60", x"00", x"E0", x"E0", x"C0", x"00", x"00", x"CE", x"80", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"08", x"1C", x"3F", x"3F", x"3F", x"3F", x"1F", x"1F", x"0F", x"0B", x"08", x"38", x"1C", x"1F", x"1F", x"1F", x"7F", x"0A", x"00", x"00", x"67", x"6D", x"7F", x"7F", x"00", x"15", x"1F", x"0F", x"05", x"02", x"14", x"74", x"3F", x"0A", x"1F", x"0F", x"0F", x"00", x"00", x"00", x"06", x"1F", x"1F", x"0F", x"0F", x"07", x"0F", x"00", x"F0", x"60", x"F0", x"F8", x"78", x"00", x"00", x"00", x"CE", x"80", x"FC", x"FE", x"7A", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"1F", x"1F", x"7F", x"30", x"00", x"00", x"07", x"0F", x"1F", x"1F", x"7F", x"0F", x"00", x"00", x"00", x"80", x"CC", x"D2", x"E0", x"20", x"00", x"00", x"00", x"80", x"4C", x"DE", x"FE", x"DE", 
															x"30", x"1F", x"0F", x"1F", x"1F", x"1F", x"1F", x"1F", x"0F", x"04", x"0C", x"0E", x"0F", x"0F", x"0F", x"07", x"20", x"F0", x"F0", x"F0", x"F8", x"FC", x"FC", x"BC", x"DE", x"4C", x"20", x"20", x"F8", x"FC", x"FC", x"BC", x"1F", x"3F", x"0F", x"0F", x"0E", x"06", x"00", x"00", x"1F", x"0F", x"0F", x"0F", x"0F", x"07", x"03", x"03", x"B8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B8", x"3C", x"00", x"C0", x"C0", x"C0", x"C0", x"80", x"07", x"0F", x"0F", x"18", x"17", x"37", x"1F", x"3F", x"07", x"0F", x"0F", x"1F", x"1F", x"3F", x"0F", x"0F", x"80", x"CC", x"D2", x"21", x"E1", x"F1", x"F2", x"F8", x"80", x"4C", x"DE", x"FF", x"DF", x"FF", x"FE", x"F8", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"7F", x"E0", x"1F", x"1F", x"1F", x"1F", x"3F", x"0F", x"07", x"0F", x"FC", x"FC", x"FE", x"1E", x"1E", x"BE", x"BC", x"00", x"FC", x"FC", x"FE", x"1E", x"1E", x"BE", x"BC", x"3E", 
															x"FE", x"14", x"00", x"40", x"EF", x"FD", x"FF", x"7F", x"01", x"2B", x"3F", x"1F", x"0B", x"12", x"34", x"64", x"80", x"00", x"00", x"8E", x"E0", x"00", x"F0", x"FE", x"60", x"C0", x"8E", x"0E", x"0E", x"FF", x"4E", x"4E", x"10", x"00", x"04", x"0F", x"1F", x"1F", x"3F", x"3F", x"0F", x"07", x"03", x"04", x"04", x"04", x"0E", x"0F", x"18", x"24", x"40", x"C0", x"C0", x"E0", x"F8", x"F8", x"F8", x"FC", x"BC", x"7C", x"7C", x"58", x"E0", x"E0", x"1F", x"07", x"2A", x"3F", x"1F", x"01", x"00", x"00", x"06", x"1F", x"BF", x"FF", x"7F", x"21", x"00", x"00", x"F0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"E0", x"F0", x"F0", x"E0", x"E0", x"C0", x"E0", x"F0", x"F0", x"E0", x"00", x"E0", x"F0", x"E0", x"00", x"00", x"CE", x"80", x"E0", x"E0", x"F8", x"F8", x"18", x"30", x"7F", x"67", x"0A", x"3F", x"3C", x"38", x"00", x"00", x"1E", x"1F", x"1F", x"3F", x"3C", x"38", x"38", x"78", 
															x"10", x"00", x"00", x"07", x"0F", x"0F", x"1F", x"1F", x"0F", x"07", x"07", x"04", x"08", x"09", x"1F", x"1F", x"10", x"00", x"40", x"DE", x"E0", x"E4", x"E0", x"FE", x"E0", x"C0", x"9E", x"DE", x"DE", x"DE", x"DE", x"DE", x"1F", x"3F", x"38", x"3C", x"1C", x"00", x"00", x"00", x"1F", x"3F", x"38", x"3C", x"1C", x"3C", x"78", x"00", x"E0", x"F0", x"78", x"38", x"78", x"00", x"00", x"00", x"FE", x"F0", x"78", x"38", x"78", x"78", x"3C", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"0F", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"F0", x"F8", x"00", x"00", x"00", x"C0", x"E0", x"D0", x"F0", x"F8", x"0B", x"08", x"08", x"00", x"00", x"37", x"7F", x"7F", x"07", x"07", x"07", x"03", x"63", x"F4", x"F8", x"FD", x"E8", x"08", x"08", x"00", x"20", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"C0", x"C0", x"C6", 
															x"7F", x"77", x"61", x"00", x"01", x"03", x"03", x"00", x"FF", x"77", x"61", x"00", x"01", x"03", x"03", x"03", x"F0", x"F9", x"F6", x"E0", x"E2", x"C0", x"80", x"00", x"CF", x"EF", x"EF", x"EF", x"EF", x"C6", x"80", x"C0", x"00", x"03", x"07", x"0F", x"0F", x"1F", x"10", x"10", x"00", x"03", x"07", x"0F", x"0F", x"1F", x"0F", x"0F", x"00", x"80", x"C0", x"E0", x"E0", x"F0", x"10", x"10", x"00", x"80", x"C0", x"A0", x"E0", x"F0", x"E0", x"E0", x"03", x"0F", x"1F", x"02", x"00", x"07", x"18", x"1F", x"03", x"03", x"00", x"05", x"07", x"02", x"43", x"42", x"F0", x"D8", x"D0", x"00", x"C0", x"80", x"2E", x"F0", x"EC", x"A0", x"2C", x"F8", x"B0", x"EE", x"EE", x"CE", x"3E", x"7F", x"7F", x"7F", x"77", x"33", x"03", x"01", x"FB", x"FE", x"FE", x"FF", x"F7", x"F3", x"43", x"01", x"80", x"F8", x"FE", x"FC", x"FC", x"F8", x"F0", x"E0", x"7F", x"26", x"22", x"C2", x"00", x"80", x"F0", x"E0", 
															x"00", x"00", x"00", x"00", x"00", x"18", x"24", x"40", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"7C", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"0F", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"0F", x"40", x"40", x"20", x"C4", x"EC", x"FE", x"FE", x"FE", x"7C", x"7C", x"3C", x"C8", x"E0", x"D2", x"FE", x"F8", x"08", x"08", x"08", x"00", x"02", x"07", x"07", x"07", x"07", x"07", x"07", x"03", x"03", x"03", x"03", x"01", x"0E", x"0E", x"0E", x"1E", x"3C", x"FC", x"F8", x"F8", x"F0", x"F0", x"F0", x"E0", x"E0", x"30", x"18", x"98", x"03", x"0F", x"0F", x"0E", x"0F", x"07", x"00", x"00", x"03", x"0F", x"0F", x"0E", x"1F", x"1F", x"0E", x"00", x"FC", x"FC", x"FE", x"18", x"18", x"08", x"00", x"00", x"FC", x"FC", x"FE", x"1E", x"1F", x"0F", x"07", x"0F", x"00", x"00", x"00", x"00", x"38", x"7C", x"FE", x"FE", x"00", x"00", x"00", x"00", x"38", x"7C", x"FA", x"FE", 
															x"18", x"10", x"10", x"03", x"07", x"0F", x"0F", x"0F", x"1F", x"0F", x"0F", x"06", x"03", x"07", x"07", x"07", x"30", x"10", x"10", x"F0", x"F8", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"10", x"F0", x"FC", x"FE", x"FE", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"0F", x"00", x"B0", x"98", x"0C", x"00", x"80", x"80", x"00", x"00", x"BE", x"9E", x"0C", x"00", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"1C", x"1C", x"1C", x"00", x"00", x"00", x"00", x"00", x"1C", x"2E", x"6F", x"FF", x"AA", x"00", x"00", x"00", x"3C", x"00", x"2A", x"00", x"3C", x"57", x"FE", x"7F", x"02", x"7F", x"55", x"7F", x"02", x"04", x"04", x"04", x"08", x"08", x"00", x"00", x"00", x"3B", x"3A", x"3B", x"34", x"34", x"1E", x"33", x"F7", x"1C", x"1C", x"1C", x"00", x"00", x"00", x"00", x"00", x"1C", x"2E", x"6F", x"FF", x"AA", x"03", x"56", x"FF", 
															x"00", x"00", x"3C", x"00", x"2A", x"00", x"3C", x"04", x"FE", x"7F", x"02", x"7F", x"55", x"7F", x"02", x"3B", x"04", x"04", x"04", x"08", x"00", x"00", x"00", x"00", x"38", x"38", x"38", x"37", x"1F", x"09", x"0D", x"3C", x"04", x"04", x"04", x"08", x"00", x"00", x"00", x"00", x"38", x"38", x"B8", x"B4", x"FC", x"C4", x"06", x"1E", x"00", x"00", x"66", x"66", x"00", x"81", x"C3", x"7E", x"00", x"3C", x"5A", x"18", x"7E", x"7E", x"3C", x"81", x"81", x"24", x"42", x"3C", x"00", x"24", x"3C", x"00", x"7E", x"DB", x"3C", x"81", x"BD", x"DB", x"42", x"3C", x"00", x"00", x"00", x"18", x"18", x"42", x"7E", x"3C", x"00", x"81", x"BD", x"E7", x"66", x"3C", x"00", x"00", x"10", x"00", x"0C", x"00", x"20", x"00", x"3C", x"00", x"0D", x"BF", x"F1", x"B9", x"9E", x"1C", x"00", x"7E", x"2A", x"00", x"3C", x"02", x"14", x"14", x"00", x"E7", x"55", x"3F", x"00", x"3C", x"7E", x"7E", x"7E", x"7E", 
															x"00", x"00", x"00", x"00", x"00", x"3C", x"00", x"3C", x"00", x"00", x"3C", x"7E", x"7E", x"42", x"FF", x"C3", x"5A", x"00", x"3C", x"00", x"24", x"00", x"3C", x"00", x"A5", x"7E", x"00", x"7E", x"5A", x"7E", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"18", x"00", x"00", x"3C", x"3C", x"3C", x"3C", x"3C", x"66", x"42", x"C3", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"5A", x"DB", x"FF", x"00", x"00", x"3C", x"00", x"24", x"00", x"3C", x"00", x"FF", x"7E", x"00", x"7E", x"5A", x"7E", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"7C", x"7C", x"DE", x"06", x"02", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"BD", x"BD", x"FF", x"42", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"7E", x"FF", x"FF", x"BD", x"BD", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7E", x"7E", x"3C", x"66", x"42", x"42", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7E", x"BD", x"FF", x"C3", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"67", x"98", x"00", x"00", x"01", x"03", x"07", x"07", x"6F", x"FF", x"FF", x"FF", x"7E", x"FF", x"FF", x"BD", x"BD", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7E", x"7E", x"7C", x"C6", x"02", x"02", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"7F", x"FF", x"AA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D7", x"FE", x"7F", x"1E", x"3F", x"3F", x"3F", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"C0", x"E0", x"F0", x"F0", x"F0", x"08", x"00", x"00", x"C0", x"E0", x"D0", x"F0", x"F8", x"F8", x"0F", x"03", x"01", x"0C", x"1E", x"1B", x"0F", x"07", x"F7", x"F7", x"F6", x"73", x"03", x"05", x"01", x"01", x"F8", x"E0", x"C0", x"00", x"38", x"F8", x"F8", x"F8", x"F0", x"70", x"30", x"E0", x"C8", x"C0", x"08", x"08", x"07", x"07", x"0F", x"0F", x"0F", x"07", x"07", x"00", x"07", x"07", x"0F", x"0F", x"0F", x"07", x"07", x"0F", x"07", x"0F", x"1F", x"1F", x"7F", x"14", x"6E", x"F7", x"07", x"0F", x"1F", x"1F", x"7F", x"0B", x"11", x"08", x"00", x"80", x"C0", x"C0", x"E0", x"00", x"C0", x"C0", x"00", x"80", x"40", x"C0", x"E0", x"C0", x"20", x"20", x"08", x"00", x"1F", x"07", x"0D", x"0F", x"1F", x"1F", x"70", x"00", x"00", x"03", x"02", x"04", x"04", x"0E", x"80", x"80", x"8E", x"E0", x"00", x"F0", x"FE", x"F0", x"60", x"4E", x"0E", x"0E", x"FF", x"4E", x"4E", x"CE", 
															x"1B", x"0F", x"0F", x"07", x"03", x"00", x"00", x"00", x"1F", x"0F", x"0F", x"07", x"03", x"00", x"01", x"00", x"E0", x"E0", x"E0", x"F0", x"E0", x"20", x"00", x"00", x"80", x"E0", x"E0", x"F8", x"F8", x"F8", x"F0", x"00", x"00", x"00", x"00", x"38", x"3C", x"1E", x"3E", x"7C", x"00", x"3E", x"7A", x"38", x"3C", x"1E", x"3E", x"7C", x"00", x"00", x"00", x"00", x"40", x"68", x"68", x"3C", x"00", x"00", x"00", x"00", x"00", x"88", x"88", x"CC", x"FE", x"F7", x"FF", x"FF", x"FF", x"FF", x"7F", x"3E", x"F8", x"5C", x"1E", x"97", x"91", x"F1", x"61", x"3E", x"5E", x"EF", x"FF", x"EF", x"CF", x"EE", x"6C", x"08", x"AE", x"1F", x"0F", x"1F", x"3D", x"1E", x"1C", x"68", x"00", x"00", x"19", x"1C", x"38", x"1D", x"1C", x"0E", x"00", x"00", x"01", x"01", x"09", x"18", x"41", x"C3", x"00", x"38", x"7C", x"3E", x"FE", x"BE", x"7E", x"6E", x"00", x"38", x"7C", x"FE", x"1A", x"4E", x"86", x"96", 
															x"6F", x"7F", x"77", x"7F", x"4F", x"0E", x"07", x"03", x"E6", x"FC", x"FC", x"7E", x"4F", x"0F", x"07", x"03", x"1C", x"9A", x"D0", x"E2", x"FF", x"FF", x"9E", x"E2", x"E4", x"66", x"28", x"60", x"C4", x"C8", x"88", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"E8", x"F8", x"F0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"00", x"00", x"10", x"20", x"30", x"1A", x"3E", x"18", x"1C", x"08", x"08", x"10", x"00", x"58", x"24", x"08", x"00", x"00", x"18", x"38", x"BA", x"7C", x"7E", x"FC", x"38", x"54", x"00", x"00", x"0C", x"3C", x"68", x"1E", x"0A", x"10", x"42", x"24", x"2E", x"BD", x"7C", x"3E", x"3E", x"51", x"F8", x"FC", x"BC", x"3C", x"1C", x"80", x"80", x"00", x"18", x"FC", x"BC", x"3E", x"1E", x"8E", x"80", x"00", x"00", x"20", x"30", x"7C", x"3C", x"28", x"18", x"00", x"49", x"B2", x"7C", x"FE", x"7D", x"7E", x"BA", x"95", 
															x"00", x"00", x"00", x"00", x"38", x"7C", x"FE", x"FE", x"00", x"00", x"00", x"00", x"38", x"7C", x"FA", x"FE", x"0F", x"10", x"1F", x"17", x"03", x"08", x"1F", x"1C", x"1F", x"1F", x"0F", x"0E", x"0C", x"07", x"03", x"03", x"E0", x"10", x"F0", x"D0", x"80", x"30", x"F0", x"F8", x"F0", x"F0", x"E0", x"E0", x"60", x"C0", x"80", x"88", x"18", x"02", x"08", x"0D", x"0E", x"07", x"07", x"00", x"07", x"07", x"0F", x"0F", x"0F", x"07", x"07", x"0F", x"78", x"38", x"B8", x"30", x"00", x"00", x"00", x"00", x"C8", x"F8", x"F8", x"F0", x"B8", x"00", x"00", x"00", x"01", x"03", x"07", x"07", x"00", x"0F", x"0B", x"0B", x"01", x"03", x"07", x"07", x"0F", x"0F", x"07", x"74", x"FC", x"FC", x"FC", x"FC", x"F0", x"60", x"00", x"00", x"F0", x"FC", x"F0", x"F0", x"F0", x"60", x"F0", x"78", x"C0", x"F8", x"FC", x"FC", x"0C", x"FC", x"EC", x"EC", x"C0", x"E0", x"C0", x"FC", x"F0", x"F0", x"70", x"10", 
															x"79", x"04", x"1F", x"17", x"7F", x"1E", x"02", x"0F", x"7E", x"7F", x"66", x"6A", x"63", x"61", x"0F", x"0F", x"CC", x"1C", x"F8", x"F8", x"F0", x"30", x"A0", x"F8", x"30", x"F0", x"30", x"30", x"F0", x"F0", x"F8", x"F8", x"0E", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"1F", x"1F", x"0F", x"00", x"00", x"00", x"00", x"38", x"38", x"78", x"78", x"78", x"70", x"00", x"00", x"38", x"38", x"78", x"78", x"78", x"70", x"70", x"38", x"C0", x"E0", x"F0", x"F0", x"00", x"F8", x"E8", x"E8", x"C0", x"E0", x"D0", x"F0", x"F8", x"F8", x"70", x"10", x"C0", x"18", x"FC", x"FC", x"FC", x"3C", x"A0", x"F8", x"30", x"E0", x"20", x"3C", x"F0", x"F0", x"F8", x"F8", x"00", x"00", x"00", x"01", x"03", x"03", x"00", x"07", x"00", x"00", x"00", x"01", x"03", x"03", x"37", x"7F", x"00", x"00", x"E0", x"F0", x"F8", x"F8", x"00", x"FC", x"00", x"00", x"E0", x"F0", x"E8", x"F8", x"FC", x"FC", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"78", x"C4", x"E4", x"78", x"86", x"86", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"35", x"00", x"0E", x"1B", x"1F", x"1F", x"1E", x"7B", x"7A", x"7B", x"73", x"35", x"11", x"1F", x"1E", x"F4", x"F4", x"E0", x"00", x"F8", x"F8", x"38", x"B8", x"B8", x"08", x"18", x"F0", x"10", x"E0", x"E0", x"E0", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"3C", x"00", x"00", x"01", x"01", x"01", x"00", x"F8", x"7C", x"70", x"F0", x"F0", x"E0", x"00", x"00", x"F8", x"60", x"70", x"F0", x"F0", x"E0", x"C0", x"E0", x"18", x"20", x"41", x"43", x"43", x"00", x"1F", x"19", x"18", x"38", x"7D", x"7F", x"7B", x"1F", x"03", x"07", x"00", x"E0", x"F0", x"F8", x"F8", x"00", x"FC", x"F4", x"00", x"E0", x"F0", x"E8", x"F8", x"FC", x"F8", x"B8", 
															x"00", x"00", x"3C", x"7E", x"7E", x"FF", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"1E", x"0F", x"0F", x"0E", x"0F", x"07", x"00", x"03", x"03", x"0F", x"0F", x"0E", x"0F", x"07", x"0E", x"E0", x"0C", x"1E", x"FE", x"1E", x"3E", x"3E", x"07", x"18", x"F8", x"F8", x"F8", x"18", x"38", x"3E", x"18", x"F0", x"E0", x"10", x"F8", x"78", x"38", x"00", x"00", x"CE", x"90", x"F0", x"F8", x"78", x"38", x"38", x"3C", x"00", x"00", x"00", x"E0", x"F0", x"F8", x"F8", x"00", x"00", x"00", x"00", x"E0", x"F0", x"E8", x"F8", x"F8", x"00", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"3C", x"3C", x"3C", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"24", x"24", x"03", x"03", x"00", x"00", x"42", x"00", x"00", x"00", x"98", x"00", x"01", x"99", x"D9", x"E0", x"78", x"2C", x"34", x"DB", x"00", x"7E", x"18", x"00", x"18", x"2C", x"34", x"18", x"00", x"00", x"00", x"3C", x"3C", x"24", x"00", x"00", x"1E", x"38", x"00", x"3C", x"18", x"3C", x"00", x"00", x"FF", x"FF", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"24", x"24", x"18", x"81", x"00", x"66", x"E7", x"5A", x"DB", x"DB", x"24", x"FF", x"66", x"00", x"00", x"3C", x"7E", x"7E", x"C3", x"81", x"81", x"42", x"18", x"7E", x"FF", x"5A", x"FF", x"DB", x"DB", x"7E", x"18", x"7E", x"FF", x"DB", x"FF", x"7E", x"7E", x"66", x"00", x"5A", x"C3", x"A5", x"81", x"81", x"42", x"66", x"66", x"FF", x"FF", x"7F", x"1E", x"14", x"16", x"33", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"3C", x"7E", x"7E", x"FF", x"7F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"77", x"55", x"55", x"55", x"55", x"77", x"00", x"00", x"77", x"55", x"55", x"55", x"55", x"77", x"00", x"00", x"01", x"03", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"03", x"01", x"01", x"01", x"01", x"00", x"00", x"07", x"01", x"07", x"04", x"04", x"07", x"00", x"00", x"07", x"01", x"07", x"04", x"04", x"07", x"00", x"00", x"02", x"06", x"0A", x"0A", x"0F", x"02", x"00", x"00", x"02", x"06", x"0A", x"0A", x"0F", x"02", x"00", x"00", x"07", x"05", x"07", x"05", x"05", x"07", x"00", x"00", x"07", x"05", x"07", x"05", x"05", x"07", x"00", x"00", x"17", x"34", x"17", x"15", x"15", x"17", x"00", x"00", x"17", x"34", x"17", x"15", x"15", x"17", x"00", x"00", x"77", x"11", x"77", x"14", x"14", x"77", x"00", x"00", x"77", x"11", x"77", x"14", x"14", x"77", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"22", x"22", x"22", x"00", x"00", x"00", x"00", x"08", x"5D", x"5D", x"5D", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5D", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"7E", x"BC", x"E6", x"43", x"03", x"07", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"7F", x"1F", x"13", x"19", x"09", x"0C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"FF", x"7E", x"FF", x"FF", x"C3", x"42", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BD", x"FF", x"FF", x"FF", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"5D", x"5D", x"5D", x"00", x"00", x"00", x"00", x"08", x"7F", x"7F", x"7F", x"5D", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"7F", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"08", x"0C", x"00", x"00", x"00", x"00", x"04", x"28", x"1C", x"0E", x"14", x"00", x"00", x"00", x"00", x"00", x"18", x"1C", x"08", x"00", x"00", x"00", x"24", x"1A", x"3C", x"3F", x"1E", x"2C", x"00", x"00", x"08", x"30", x"20", x"50", x"38", x"10", x"00", x"3A", x"7C", x"7C", x"F8", x"FA", x"FE", x"7C", x"38", x"00", x"00", x"28", x"30", x"60", x"24", x"10", x"00", x"18", x"BC", x"7D", x"FE", x"FB", x"FC", x"7C", x"3A", 
															x"1C", x"3A", x"3A", x"7F", x"7F", x"3E", x"3E", x"1C", x"3C", x"7E", x"7E", x"7F", x"7F", x"7E", x"7E", x"3C", x"04", x"0A", x"1A", x"1E", x"1E", x"1E", x"0E", x"04", x"1C", x"3E", x"3E", x"3E", x"3E", x"3E", x"3E", x"1C", x"00", x"14", x"0C", x"0C", x"0C", x"0C", x"04", x"00", x"18", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"18", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"10", x"92", x"44", x"00", x"44", x"82", x"10", x"10", x"10", x"92", x"44", x"00", x"44", x"82", x"10", x"10", x"3F", x"3E", x"3F", x"3E", x"3C", x"1E", x"33", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"7F", x"FF", x"AA", x"03", x"56", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"7F", x"3E", x"7F", x"7F", x"7F", x"3E", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3C", x"3C", x"3C", x"3F", x"1F", x"09", x"0D", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"7E", x"BD", x"BD", x"FF", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"BC", x"BC", x"FC", x"C4", x"06", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"81", x"BD", x"FF", x"7E", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1D", x"BF", x"F9", x"B9", x"BC", x"1C", x"1C", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"3F", x"3C", x"3E", x"6A", x"6A", x"7A", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"7E", x"3C", x"7E", x"7E", x"7E", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"3C", x"3C", x"3C", x"66", x"42", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"7C", x"7C", x"DE", x"02", x"02", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"BD", x"BD", x"FF", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"7F", x"00", x"00", x"00", x"00", x"00", x"1C", x"3A", x"7F", x"03", x"0F", x"03", x"0E", x"1D", x"00", x"18", x"1D", x"03", x"0F", x"00", x"01", x"02", x"0F", x"40", x"40", x"F8", x"FC", x"80", x"D8", x"F8", x"30", x"3E", x"F0", x"F8", x"FC", x"78", x"24", x"04", x"0E", x"0E", x"0E", x"3E", x"7F", x"7F", x"7F", x"77", x"33", x"03", x"01", x"FB", x"FE", x"FE", x"FF", x"F7", x"F3", x"43", x"01", 
															x"80", x"F8", x"FE", x"FC", x"FC", x"F8", x"F0", x"E0", x"7F", x"26", x"22", x"C2", x"00", x"80", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"3E", x"3E", x"73", x"40", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"FC", x"7C", x"F8", x"00", x"00", x"3C", x"7E", x"7E", x"FF", x"0F", x"4F", x"F8", x"F8", x"F8", x"F0", x"07", x"07", x"03", x"02", x"4F", x"0F", x"1F", x"FF", x"7F", x"FD", x"FD", x"FD", x"03", x"07", x"03", x"1E", x"14", x"16", x"33", x"F7", x"FC", x"F9", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"7C", x"F8", x"F8", x"00", x"3C", x"7E", x"7E", x"FF", x"0F", x"4F", x"4F", x"F8", x"F8", x"F0", x"07", x"07", x"03", x"12", x"36", x"0F", x"1F", x"FF", x"7F", x"FD", x"FD", x"ED", x"C9", 
															x"7F", x"7B", x"1F", x"3F", x"3C", x"38", x"00", x"00", x"1E", x"1F", x"1F", x"3F", x"3C", x"38", x"38", x"78", x"F0", x"F0", x"F0", x"F8", x"78", x"38", x"00", x"00", x"CE", x"90", x"F0", x"F8", x"78", x"38", x"38", x"3C", x"3C", x"98", x"BC", x"E6", x"42", x"03", x"03", x"0E", x"C2", x"76", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F8", x"F0", x"07", x"07", x"53", x"7E", x"70", x"0F", x"1F", x"FF", x"7F", x"FD", x"AD", x"81", x"AF", x"00", x"00", x"1E", x"13", x"19", x"09", x"0C", x"3C", x"7F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"FF", x"FF", x"FF", x"FF", x"E7", x"00", x"3C", x"7E", x"C3", x"A5", x"81", x"BD", x"FF", x"FF", x"81", x"E7", x"66", x"66", x"81", x"81", x"C3", x"42", x"FF", x"18", x"18", x"5A", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", 
															x"00", x"81", x"81", x"C3", x"42", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"3C", x"3C", x"7E", x"3C", x"00", x"00", x"00", x"00", x"0C", x"04", x"04", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"C3", x"C3", x"81", x"81", x"00", x"FF", x"FF", x"7E", x"FF", x"7E", x"7E", x"7E", x"FF", x"00", x"00", x"00", x"3C", x"66", x"42", x"42", x"C3", x"FF", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"81", x"FF", x"81", x"81", x"00", x"00", x"FF", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"FF", x"FF", x"FF", x"00", x"00", x"3C", x"7E", x"7E", x"81", x"A5", x"FF", x"00", x"00", x"00", x"C3", x"C3", x"81", x"81", x"00", x"FF", x"FF", x"7E", x"FF", x"7E", x"7E", x"7E", x"FF", x"00", x"00", x"00", x"7C", x"C6", x"02", x"02", x"03", x"FF", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"02", x"42", x"43", x"C1", x"C0", x"03", x"C3", x"00", x"18", x"3C", x"3C", x"3E", x"38", x"7E", x"7C", x"C0", x"7E", x"FF", x"FF", x"FF", x"7F", x"7F", x"3E", x"3F", x"7F", x"C3", x"81", x"D5", x"D5", x"E3", x"7E", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"7F", x"40", x"40", x"40", x"40", x"40", x"40", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"66", x"66", x"66", x"00", x"00", x"00", x"00", x"00", x"66", x"22", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"82", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"82", x"FE", x"1C", x"3E", x"FF", x"38", x"6D", x"DF", x"0F", x"3C", x"1C", x"3A", x"FF", x"07", x"12", x"20", x"70", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"02", x"02", x"02", x"02", x"02", x"02", x"FE", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"C4", x"E4", x"78", x"86", x"86", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"06", x"06", x"06", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"DE", x"CC", x"7A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"7C", x"38", x"7C", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"0E", x"1C", x"38", x"70", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"10", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"20", x"20", x"00", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6C", x"FE", x"FE", x"FE", x"7C", x"38", x"10", x"70", x"70", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"60", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"70", x"70", x"00", x"00", x"00", x"00", x"00", x"C0", x"40", x"60", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", 
															x"00", x"FF", x"60", x"6F", x"6F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"06", x"E6", x"E6", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"3F", x"20", x"20", x"20", x"3F", x"20", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"FC", x"04", x"04", x"04", x"FC", x"04", x"04", x"00", x"01", x"01", x"03", x"FF", x"00", x"10", x"10", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"03", x"7F", x"01", x"21", x"21", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"30", x"F7", x"00", x"01", x"01", x"03", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"63", x"EF", x"01", x"01", x"01", x"03", x"7F", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"10", x"10", x"30", x"F7", x"00", x"01", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"21", x"21", x"63", x"EF", x"01", x"01", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"A0", x"A0", x"AA", x"AA", x"AA", x"AA", x"AA", x"00", x"7F", x"7F", x"75", x"7F", x"7F", x"7F", x"7F", x"00", x"0B", x"0B", x"AB", x"AB", x"AB", x"AB", x"AB", x"00", x"FD", x"FD", x"5D", x"FD", x"FD", x"FD", x"FD", x"A0", x"A0", x"A0", x"A0", x"A0", x"A0", x"A0", x"A0", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"00", x"00", x"00", x"30", x"3F", x"1F", x"00", x"30", x"00", x"FF", x"FF", x"CF", x"E0", x"FF", x"FF", x"CF", x"00", x"01", x"01", x"19", x"F9", x"F1", x"01", x"19", x"00", x"FF", x"FF", x"E7", x"0F", x"FF", x"FF", x"E7", 
															x"3F", x"1F", x"00", x"30", x"3F", x"1F", x"00", x"30", x"E0", x"FF", x"FF", x"CF", x"E0", x"FF", x"FF", x"CF", x"F9", x"F1", x"01", x"19", x"F9", x"F1", x"01", x"19", x"0F", x"FF", x"FF", x"E7", x"0F", x"FF", x"FF", x"E7", x"3F", x"1F", x"00", x"30", x"3F", x"1F", x"00", x"00", x"E0", x"FF", x"FF", x"CF", x"E0", x"FF", x"FF", x"FF", x"F9", x"F1", x"01", x"19", x"F9", x"F1", x"01", x"01", x"0F", x"FF", x"FF", x"E7", x"0F", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"1F", x"3F", x"3C", x"35", x"35", x"00", x"FF", x"C0", x"80", x"80", x"80", x"A8", x"E0", x"00", x"00", x"00", x"70", x"78", x"78", x"D8", x"D8", x"00", x"FE", x"06", x"02", x"02", x"02", x"2A", x"0E", x"3D", x"3C", x"3F", x"3F", x"3F", x"34", x"35", x"3D", x"E0", x"A0", x"80", x"80", x"80", x"88", x"80", x"80", x"F8", x"78", x"78", x"78", x"78", x"58", x"D8", x"F8", x"0E", x"0A", x"02", x"02", x"02", x"22", x"02", x"02", 
															x"3D", x"3C", x"3F", x"3F", x"37", x"34", x"3D", x"3D", x"80", x"80", x"A0", x"E0", x"E8", x"A0", x"80", x"80", x"F8", x"78", x"78", x"78", x"58", x"58", x"F8", x"F8", x"02", x"02", x"0A", x"0E", x"2E", x"0A", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"07", x"00", x"01", x"00", x"00", x"01", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"00", x"00", x"80", x"80", x"00", x"80", x"00", x"C0", x"0F", x"0F", x"1F", x"1F", x"1F", x"1F", x"0F", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"1F", x"0F", x"0F", x"60", x"20", x"B0", x"F0", x"F0", x"F0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"07", x"00", x"3F", x"3F", x"74", x"74", x"E4", x"FF", x"07", x"00", x"00", x"1B", x"10", x"30", x"20", x"00", x"C0", x"00", x"F8", x"F8", x"5C", x"5C", x"4E", x"FE", x"C0", x"00", x"00", x"B0", x"10", x"18", x"08", x"00", 
															x"00", x"00", x"0F", x"1F", x"3F", x"00", x"1F", x"00", x"00", x"00", x"0F", x"10", x"3F", x"1F", x"00", x"00", x"00", x"00", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"09", x"09", x"09", x"09", x"00", x"7F", x"FC", x"F8", x"FF", x"FF", x"00", x"FF", x"00", x"7F", x"FC", x"FB", x"00", x"FF", x"FF", x"00", x"00", x"03", x"05", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"24", x"24", x"24", x"24", x"00", x"FF", x"3C", x"18", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"3C", x"DB", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"81", x"81", x"BD", x"00", x"00", x"FF", x"00", x"FF", x"81", x"81", x"BD", x"00", x"FF", x"FE", x"00", x"FD", x"81", x"83", x"B3", x"07", x"00", x"FE", x"00", x"FC", x"80", x"81", x"B1", x"03", x"E6", x"2F", x"0C", x"FF", x"FF", x"00", x"FF", x"00", x"E3", x"27", x"C7", x"0F", x"FF", x"FF", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"1F", x"60", x"FF", x"C0", x"FF", x"8C", x"F9", x"12", x"F4", x"3F", x"7F", x"7F", x"FF", x"FF", x"FE", x"FC", x"F8", x"24", x"E8", x"48", x"D0", x"90", x"20", x"E0", x"00", x"F8", x"F0", x"F0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F8", x"06", x"FF", x"03", x"FF", x"31", x"9F", x"48", x"2F", x"FC", x"FE", x"FE", x"FF", x"FF", x"7F", x"3F", x"1F", x"24", x"17", x"12", x"0B", x"09", x"04", x"07", x"00", x"1F", x"0F", x"0F", x"07", x"07", x"03", x"00", x"00", 
															x"00", x"01", x"01", x"03", x"FF", x"08", x"14", x"15", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"13", x"7F", x"01", x"61", x"A1", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"32", x"F7", x"04", x"05", x"09", x"0B", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"63", x"EF", x"81", x"61", x"11", x"03", x"7F", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"10", x"10", x"30", x"F7", x"00", x"01", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"21", x"21", x"63", x"EF", x"01", x"01", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"21", x"21", x"13", x"FF", x"08", x"14", x"15", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"29", x"51", x"13", x"7F", x"01", x"69", x"A5", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"32", x"F7", x"04", x"15", x"29", x"4B", x"FF", x"14", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"63", x"EF", x"81", x"69", x"11", x"23", x"7F", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"12", x"12", x"34", x"F7", x"00", x"01", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"29", x"A1", x"63", x"EF", x"01", x"01", x"01", x"03", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"62", x"10", x"00", x"09", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"84", x"A0", x"C0", x"4C", x"04", x"60", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"40", x"12", x"04", x"0F", x"2E", x"64", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"68", x"4C", x"18", x"14", x"40", x"48", x"DC", x"80", 
															x"00", x"00", x"00", x"FF", x"01", x"01", x"01", x"03", x"46", x"14", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"01", x"01", x"01", x"01", x"18", x"B0", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"30", x"16", x"00", x"24", x"33", x"76", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"D0", x"D4", x"84", x"2C", x"04", x"20", x"74", x"00", x"00", x"00", x"FF", x"01", x"01", x"01", x"03", x"41", x"63", x"08", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"01", x"01", x"01", x"01", x"10", x"44", x"0C", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"20", x"72", x"14", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"80", x"6C", x"C4", x"00", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"20", x"72", x"04", x"30", x"3F", x"1F", x"00", x"00", x"00", x"00", x"00", x"40", x"E0", x"FF", x"FF", x"FF", x"0C", x"64", x"C0", x"18", x"F9", x"F1", x"01", x"01", x"00", x"00", x"00", x"04", x"0F", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"30", x"3F", x"1F", x"00", x"00", x"00", x"00", x"00", x"40", x"E0", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"18", x"F9", x"F1", x"01", x"01", x"00", x"00", x"00", x"04", x"0F", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"30", x"A1", x"A0", x"A0", x"A0", x"20", x"75", x"02", x"08", x"7C", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"08", x"9B", x"0B", x"0B", x"0B", x"30", x"66", x"02", x"00", x"6D", x"FD", x"FD", x"FD", 
															x"00", x"00", x"00", x"30", x"A1", x"A0", x"A0", x"A0", x"00", x"00", x"00", x"08", x"7C", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"08", x"9B", x"0B", x"0B", x"0B", x"00", x"00", x"00", x"00", x"6D", x"FD", x"FD", x"FD", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"62", x"4C", x"01", x"33", x"15", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"4C", x"40", x"20", x"08", x"98", x"80", x"00", x"00", x"00", x"00", x"03", x"03", x"01", x"0D", x"1D", x"00", x"00", x"00", x"00", x"00", x"01", x"0D", x"1D", x"00", x"00", x"00", x"00", x"80", x"C0", x"60", x"20", x"00", x"00", x"00", x"80", x"00", x"C0", x"E0", x"E0", x"1B", x"19", x"1C", x"08", x"04", x"1C", x"0E", x"0F", x"1B", x"19", x"1C", x"08", x"04", x"1C", x"0E", x"0F", x"B0", x"F0", x"A0", x"00", x"D0", x"70", x"E0", x"60", x"F0", x"F0", x"A0", x"00", x"D0", x"70", x"E0", x"60", 
															x"00", x"00", x"03", x"0B", x"18", x"12", x"32", x"38", x"00", x"00", x"00", x"08", x"18", x"12", x"32", x"38", x"00", x"00", x"00", x"80", x"30", x"58", x"48", x"6C", x"00", x"00", x"80", x"00", x"30", x"78", x"78", x"7C", x"10", x"00", x"00", x"04", x"30", x"18", x"1C", x"0E", x"10", x"00", x"00", x"04", x"30", x"18", x"1C", x"0E", x"38", x"24", x"00", x"18", x"50", x"30", x"60", x"00", x"38", x"24", x"00", x"18", x"50", x"30", x"60", x"00", x"00", x"00", x"3F", x"3F", x"74", x"74", x"E4", x"FF", x"00", x"00", x"00", x"1B", x"10", x"30", x"20", x"00", x"00", x"00", x"F8", x"F8", x"5C", x"5C", x"4E", x"FE", x"00", x"00", x"00", x"B0", x"10", x"18", x"08", x"00", x"00", x"02", x"37", x"60", x"40", x"E0", x"50", x"00", x"00", x"01", x"30", x"60", x"40", x"E0", x"50", x"00", x"00", x"00", x"00", x"32", x"A8", x"90", x"06", x"04", x"00", x"00", x"00", x"32", x"B8", x"90", x"06", x"0C", 
															x"20", x"00", x"28", x"70", x"60", x"3A", x"30", x"18", x"20", x"00", x"28", x"70", x"60", x"3A", x"30", x"18", x"19", x"12", x"00", x"26", x"24", x"0C", x"18", x"00", x"19", x"12", x"00", x"26", x"24", x"0C", x"18", x"00", x"00", x"22", x"60", x"D0", x"80", x"80", x"00", x"00", x"00", x"20", x"60", x"D0", x"80", x"80", x"00", x"00", x"00", x"02", x"05", x"03", x"00", x"08", x"01", x"00", x"00", x"02", x"07", x"03", x"08", x"08", x"01", x"00", x"00", x"00", x"20", x"00", x"80", x"C0", x"C0", x"60", x"00", x"00", x"20", x"00", x"80", x"C0", x"C0", x"60", x"00", x"00", x"00", x"00", x"01", x"05", x"03", x"0E", x"00", x"00", x"00", x"00", x"01", x"05", x"03", x"0E", x"00", x"00", x"00", x"30", x"38", x"3C", x"34", x"34", x"00", x"FF", x"C0", x"80", x"80", x"80", x"A8", x"E0", x"00", x"00", x"00", x"18", x"38", x"78", x"58", x"58", x"00", x"FE", x"06", x"02", x"02", x"02", x"2A", x"0E", 
															x"38", x"38", x"38", x"38", x"3C", x"34", x"34", x"3C", x"A0", x"A0", x"80", x"80", x"80", x"88", x"80", x"80", x"38", x"38", x"38", x"38", x"78", x"58", x"58", x"78", x"0A", x"0A", x"02", x"02", x"02", x"22", x"02", x"02", x"38", x"38", x"38", x"38", x"34", x"34", x"38", x"30", x"80", x"80", x"A0", x"E0", x"E8", x"A0", x"80", x"80", x"38", x"38", x"38", x"38", x"58", x"58", x"38", x"18", x"02", x"02", x"0A", x"0E", x"2E", x"0A", x"02", x"02", x"00", x"00", x"00", x"00", x"60", x"70", x"70", x"70", x"00", x"FF", x"C0", x"80", x"80", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"0C", x"1C", x"1C", x"1C", x"00", x"FE", x"06", x"02", x"02", x"02", x"06", x"06", x"70", x"70", x"70", x"70", x"70", x"70", x"70", x"70", x"C0", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"06", x"06", x"02", x"02", x"02", x"02", x"02", x"02", 
															x"70", x"70", x"70", x"70", x"70", x"70", x"70", x"60", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"0C", x"02", x"02", x"06", x"06", x"06", x"06", x"02", x"02", x"00", x"00", x"00", x"00", x"40", x"40", x"40", x"40", x"00", x"FF", x"C0", x"80", x"80", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"04", x"04", x"04", x"04", x"00", x"FE", x"06", x"02", x"02", x"02", x"06", x"06", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"C0", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"06", x"06", x"02", x"02", x"02", x"02", x"02", x"02", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"02", x"02", x"06", x"06", x"06", x"06", x"02", x"02", 
															x"7F", x"18", x"1F", x"0F", x"06", x"04", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"30", x"F0", x"E0", x"C0", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"06", x"07", x"07", x"07", x"07", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"04", x"04", x"04", x"04", x"06", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"2C", x"02", x"00", x"20", x"74", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"10", x"4A", x"C2", x"16", 
															x"FF", x"7F", x"00", x"BF", x"81", x"C1", x"CD", x"E0", x"00", x"7F", x"00", x"3F", x"01", x"81", x"8D", x"C0", x"67", x"F4", x"30", x"FF", x"FF", x"00", x"FF", x"00", x"C7", x"E4", x"E3", x"F0", x"FF", x"FF", x"00", x"00", x"C0", x"A0", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"90", x"90", x"90", x"90", x"00", x"FE", x"3F", x"1F", x"FF", x"FF", x"00", x"FF", x"00", x"FE", x"3F", x"DF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"F0", x"F8", x"FC", x"00", x"F0", x"00", x"00", x"00", x"F0", x"08", x"FC", x"F0", x"00", x"00", x"1E", x"0E", x"0A", x"CA", x"CA", x"4A", x"4E", x"4E", x"00", x"00", x"00", x"C0", x"C0", x"40", x"40", x"40", x"4E", x"4E", x"4A", x"4A", x"4A", x"4A", x"4E", x"4E", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", 
															x"00", x"00", x"00", x"FF", x"00", x"11", x"AA", x"44", x"00", x"00", x"00", x"FF", x"00", x"11", x"AA", x"44", x"78", x"70", x"50", x"53", x"53", x"52", x"72", x"72", x"00", x"00", x"00", x"03", x"03", x"02", x"02", x"02", x"72", x"72", x"52", x"52", x"52", x"52", x"72", x"72", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"FF", x"00", x"88", x"55", x"22", x"00", x"00", x"00", x"FF", x"00", x"88", x"55", x"22", x"FF", x"FF", x"E0", x"C0", x"CF", x"CC", x"C9", x"CB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"01", x"00", x"FE", x"06", x"F2", x"FA", x"00", x"00", x"02", x"01", x"01", x"09", x"05", x"05", x"CB", x"CB", x"CB", x"CB", x"C9", x"CC", x"EF", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"FA", x"FA", x"FA", x"FA", x"F2", x"06", x"FC", x"01", x"05", x"05", x"05", x"05", x"0D", x"F9", x"03", x"FE", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"00", x"00", x"00", x"00", x"7F", x"7F", x"1F", x"1B", x"00", x"00", x"00", x"00", x"08", x"08", x"F8", x"E8", x"00", x"00", x"00", x"00", x"F6", x"F6", x"F8", x"F8", x"1F", x"1F", x"3F", x"00", x"3F", x"1F", x"1F", x"1F", x"17", x"1B", x"37", x"00", x"3B", x"17", x"1B", x"17", x"E8", x"E8", x"F4", x"00", x"EC", x"E8", x"E8", x"E8", x"F8", x"F8", x"FC", x"00", x"FC", x"F8", x"F8", x"F8", x"1F", x"1F", x"3F", x"00", x"3F", x"1F", x"1F", x"1F", x"1B", x"17", x"3B", x"00", x"37", x"1B", x"17", x"1B", x"E8", x"E8", x"F4", x"00", x"EC", x"E8", x"E8", x"E8", x"F8", x"F8", x"FC", x"00", x"FC", x"F8", x"F8", x"F8", x"1F", x"00", x"00", x"00", x"70", x"38", x"FF", x"00", x"1F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"F8", x"08", x"08", x"00", x"0E", x"1C", x"FF", x"00", x"F8", x"F6", x"F6", x"00", x"00", x"00", x"00", x"00", 
															x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"F8", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"F8", x"F6", x"F6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0F", x"1F", x"1F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"C0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"0F", x"1F", x"1F", x"1F", x"1F", x"1D", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"E0", x"E0", x"C0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"00", x"08", x"08", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"C0", x"00", x"40", x"40", x"C0", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"EF", x"EF", x"CF", x"0A", x"FE", x"FE", x"FE", x"00", x"EF", x"E0", x"CD", x"08", x"FC", x"FC", x"FE", x"00", x"EF", x"FF", x"EF", x"2A", x"FE", x"FE", x"FE", x"00", x"EF", x"49", x"C5", x"00", x"D4", x"D4", x"FE", x"AF", x"17", x"AE", x"44", x"AE", x"17", x"AF", x"40", x"A8", x"10", x"A9", x"43", x"A9", x"10", x"A8", x"40", x"FF", x"7B", x"FD", x"00", x"FD", x"7B", x"FF", x"00", x"00", x"84", x"02", x"FF", x"02", x"84", x"00", x"00", x"AA", x"91", x"AA", x"84", x"AA", x"91", x"AA", x"04", x"2A", x"11", x"2A", x"04", x"2A", x"11", x"2A", x"04", x"AA", x"11", x"AA", x"44", x"AA", x"11", x"AA", x"44", x"AA", x"11", x"AA", x"44", x"AA", x"11", x"AA", x"44", 
															x"D5", x"C8", x"D5", x"42", x"D5", x"C8", x"D5", x"02", x"15", x"08", x"15", x"82", x"15", x"08", x"15", x"02", x"FF", x"BD", x"7E", x"00", x"7E", x"BD", x"FF", x"00", x"00", x"42", x"81", x"FF", x"81", x"42", x"00", x"00", x"57", x"8B", x"57", x"22", x"57", x"8B", x"57", x"20", x"54", x"88", x"54", x"21", x"54", x"88", x"54", x"20", x"55", x"88", x"55", x"22", x"55", x"88", x"55", x"22", x"55", x"88", x"55", x"22", x"55", x"88", x"55", x"22", x"00", x"E0", x"5F", x"60", x"60", x"5F", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"FA", x"06", x"06", x"FA", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"0E", x"0E", x"07", x"07", x"03", x"00", x"00", x"00", x"06", x"02", x"03", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"46", x"6E", x"56", x"56", x"46", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"2C", x"46", x"46", x"7E", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"46", x"46", x"7C", x"48", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"18", x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"46", x"46", x"46", x"46", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"30", x"30", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"46", x"46", x"46", x"46", x"46", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"46", x"40", x"4E", x"46", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"60", x"60", x"60", x"60", x"60", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"07", x"0E", x"0E", x"00", x"00", x"00", x"00", x"00", x"03", x"02", x"06", x"FC", x"EF", x"EF", x"CF", x"FC", x"FE", x"FE", x"FE", x"00", x"29", x"29", x"09", x"00", x"3E", x"3E", x"FE", x"C6", x"EF", x"EF", x"FF", x"CE", x"FE", x"FE", x"FE", x"00", x"29", x"29", x"01", x"08", x"38", x"38", x"FE", x"78", x"EF", x"EF", x"CF", x"FE", x"FE", x"FE", x"FE", x"40", x"83", x"29", x"09", x"00", x"38", x"38", x"FE", x"78", x"EF", x"EF", x"FF", x"0E", x"FE", x"FE", x"FE", x"00", x"23", x"2F", x"83", x"08", x"38", x"82", x"FE", x"FE", x"EF", x"EF", x"FF", x"C8", x"FE", x"FE", x"FE", x"00", x"2F", x"2F", x"03", x"08", x"3E", x"00", x"FE", 
															x"40", x"EF", x"EF", x"CF", x"08", x"FE", x"FE", x"FE", x"40", x"EF", x"EF", x"CF", x"08", x"FE", x"FE", x"FE", x"00", x"EF", x"EF", x"CF", x"08", x"FE", x"FE", x"FE", x"00", x"EF", x"EF", x"CF", x"08", x"FE", x"FE", x"FE", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"F8", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"7C", x"7C", x"7C", x"7C", x"7C", x"7C", x"7C", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7C", x"7C", x"7C", x"7C", x"7C", x"7C", x"7C", x"7C", x"C0", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"F3", x"F9", x"F8", x"FC", x"FC", x"FC", x"FC", 
															x"5F", x"F0", x"C0", x"C0", x"80", x"80", x"80", x"80", x"40", x"8F", x"BF", x"3F", x"7F", x"7F", x"7F", x"7F", x"80", x"80", x"00", x"00", x"00", x"80", x"C0", x"E0", x"7F", x"7F", x"7F", x"7F", x"3F", x"BF", x"DF", x"E7", x"00", x"00", x"00", x"00", x"00", x"02", x"06", x"1E", x"FC", x"FC", x"FC", x"F8", x"F8", x"F2", x"C6", x"1E", x"80", x"80", x"80", x"80", x"08", x"FE", x"FE", x"FE", x"7C", x"7C", x"7C", x"7C", x"08", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"10", x"18", x"3C", x"FF", x"FF", x"EF", x"EF", x"C7", x"D7", x"9B", x"3D", x"00", x"01", x"03", x"0F", x"03", x"00", x"00", x"00", x"FC", x"F9", x"E3", x"8F", x"E3", x"F8", x"FC", x"FC", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC");

	constant TEST2_CHR_ROM : CHR_ROM_ARRAY := (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"00",x"6C",x"6C",x"6C",x"00",x"00",x"00",x"00",x"00",x"6C",x"6C",x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"6C",x"FE",x"6C",x"6C",x"FE",x"6C",x"00",x"00",x"6C",x"FE",x"6C",x"6C",x"FE",x"6C",x"00",
															x"18",x"3E",x"60",x"3C",x"06",x"7C",x"18",x"00",x"18",x"3E",x"60",x"3C",x"06",x"7C",x"18",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"46",x"00",x"62",x"66",x"0C",x"18",x"30",x"66",x"46",x"00",x"1C",x"36",x"1C",x"38",x"6B",x"66",x"3B",x"00",x"1C",x"36",x"1C",x"38",x"6B",x"66",x"3B",x"00",x"0C",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",x"0C",x"0C",x"0C",x"00",x"00",x"00",x"00",x"00",
															x"06",x"0C",x"18",x"18",x"18",x"0C",x"06",x"00",x"06",x"0C",x"18",x"18",x"18",x"0C",x"06",x"00",x"60",x"30",x"18",x"18",x"18",x"30",x"60",x"00",x"60",x"30",x"18",x"18",x"18",x"30",x"60",x"00",x"00",x"66",x"3C",x"FF",x"3C",x"66",x"00",x"00",x"00",x"66",x"3C",x"FF",x"3C",x"66",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",
															x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"60",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"60",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"60",x"00",x"02",x"06",x"0C",x"18",x"30",x"60",x"40",x"00",x"02",x"06",x"0C",x"18",x"30",x"60",x"40",x"00",
															x"38",x"4C",x"CE",x"C6",x"E6",x"64",x"38",x"00",x"38",x"4C",x"CE",x"C6",x"E6",x"64",x"38",x"00",x"18",x"38",x"18",x"18",x"18",x"18",x"7E",x"00",x"18",x"38",x"18",x"18",x"18",x"18",x"7E",x"00",x"7C",x"C6",x"0E",x"3C",x"78",x"E0",x"FE",x"00",x"7C",x"C6",x"0E",x"3C",x"78",x"E0",x"FE",x"00",x"7E",x"0C",x"18",x"3C",x"06",x"C6",x"7C",x"00",x"7E",x"0C",x"18",x"3C",x"06",x"C6",x"7C",x"00",
															x"1C",x"3C",x"6C",x"CC",x"FE",x"0C",x"0C",x"00",x"1C",x"3C",x"6C",x"CC",x"FE",x"0C",x"0C",x"00",x"FC",x"C0",x"FC",x"06",x"06",x"C6",x"7C",x"00",x"FC",x"C0",x"FC",x"06",x"06",x"C6",x"7C",x"00",x"3C",x"60",x"C0",x"FC",x"C6",x"C6",x"7C",x"00",x"3C",x"60",x"C0",x"FC",x"C6",x"C6",x"7C",x"00",x"FE",x"C6",x"0C",x"18",x"30",x"30",x"30",x"00",x"FE",x"C6",x"0C",x"18",x"30",x"30",x"30",x"00",
															x"78",x"C4",x"E4",x"78",x"86",x"86",x"7C",x"00",x"78",x"C4",x"E4",x"78",x"86",x"86",x"7C",x"00",x"7C",x"C6",x"C6",x"7E",x"06",x"0C",x"78",x"00",x"7C",x"C6",x"C6",x"7E",x"06",x"0C",x"78",x"00",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"60",x"00",x"18",x"18",x"00",x"00",x"18",x"18",x"60",
															x"00",x"18",x"30",x"60",x"30",x"18",x"00",x"00",x"00",x"18",x"30",x"60",x"30",x"18",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"7E",x"00",x"00",x"00",x"18",x"0C",x"06",x"0C",x"18",x"00",x"00",x"00",x"18",x"0C",x"06",x"0C",x"18",x"00",x"00",x"7C",x"C6",x"06",x"1C",x"30",x"00",x"30",x"00",x"7C",x"C6",x"06",x"1C",x"30",x"00",x"30",x"00",
															x"3C",x"66",x"6E",x"6A",x"6E",x"60",x"3E",x"00",x"3C",x"66",x"6E",x"6A",x"6E",x"60",x"3E",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"38",x"6C",x"C6",x"C6",x"FE",x"C6",x"C6",x"00",x"FC",x"C6",x"C6",x"FC",x"C6",x"C6",x"FC",x"00",x"FC",x"C6",x"C6",x"FC",x"C6",x"C6",x"FC",x"00",x"3C",x"66",x"C0",x"C0",x"C0",x"66",x"3C",x"00",x"3C",x"66",x"C0",x"C0",x"C0",x"66",x"3C",x"00",
															x"F8",x"CC",x"C6",x"C6",x"C6",x"CC",x"F8",x"00",x"F8",x"CC",x"C6",x"C6",x"C6",x"CC",x"F8",x"00",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"FE",x"00",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"FE",x"00",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"C0",x"00",x"FE",x"C0",x"C0",x"FC",x"C0",x"C0",x"C0",x"00",x"3E",x"60",x"C0",x"CE",x"C6",x"66",x"3E",x"00",x"3E",x"60",x"C0",x"CE",x"C6",x"66",x"3E",x"00",
															x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"00",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"1E",x"06",x"06",x"06",x"C6",x"C6",x"7C",x"00",x"1E",x"06",x"06",x"06",x"C6",x"C6",x"7C",x"00",x"C6",x"CC",x"D8",x"F0",x"D8",x"CC",x"C6",x"00",x"C6",x"CC",x"D8",x"F0",x"D8",x"CC",x"C6",x"00",
															x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00",x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"00",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"00",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"00",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",
															x"FC",x"C6",x"C6",x"FC",x"C0",x"C0",x"C0",x"00",x"FC",x"C6",x"C6",x"FC",x"C0",x"C0",x"C0",x"00",x"7C",x"C6",x"C6",x"C6",x"DA",x"CC",x"76",x"00",x"7C",x"C6",x"C6",x"C6",x"DA",x"CC",x"76",x"00",x"FC",x"C6",x"C6",x"FC",x"D8",x"CC",x"C6",x"00",x"FC",x"C6",x"C6",x"FC",x"D8",x"CC",x"C6",x"00",x"7C",x"C6",x"C0",x"7C",x"06",x"C6",x"7C",x"00",x"7C",x"C6",x"C0",x"7C",x"06",x"C6",x"7C",x"00",
															x"FC",x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"FC",x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"C6",x"C6",x"C6",x"EE",x"7C",x"38",x"10",x"00",x"C6",x"C6",x"C6",x"EE",x"7C",x"38",x"10",x"00",x"C6",x"C6",x"D6",x"FE",x"FE",x"EE",x"C6",x"00",x"C6",x"C6",x"D6",x"FE",x"FE",x"EE",x"C6",x"00",
															x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"C6",x"EE",x"7C",x"38",x"7C",x"EE",x"C6",x"00",x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"00",x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"00",x"FE",x"0E",x"1C",x"38",x"70",x"E0",x"FE",x"00",x"FE",x"0E",x"1C",x"38",x"70",x"E0",x"FE",x"00",x"1E",x"18",x"18",x"18",x"18",x"18",x"1E",x"00",x"1E",x"18",x"18",x"18",x"18",x"18",x"1E",x"00",
															x"40",x"60",x"30",x"18",x"0C",x"06",x"02",x"00",x"40",x"60",x"30",x"18",x"0C",x"06",x"02",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"10",x"38",x"6C",x"C6",x"00",x"00",x"00",x"00",x"10",x"38",x"6C",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",
															x"C0",x"60",x"30",x"00",x"00",x"00",x"00",x"00",x"C0",x"60",x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"0C",x"7C",x"CC",x"76",x"00",x"00",x"00",x"78",x"0C",x"7C",x"CC",x"76",x"00",x"C0",x"C0",x"F8",x"CC",x"CC",x"CC",x"F8",x"00",x"C0",x"C0",x"F8",x"CC",x"CC",x"CC",x"F8",x"00",x"00",x"00",x"78",x"CC",x"C0",x"CC",x"78",x"00",x"00",x"00",x"78",x"CC",x"C0",x"CC",x"78",x"00",
															x"0C",x"0C",x"7C",x"CC",x"CC",x"CC",x"7C",x"00",x"0C",x"0C",x"7C",x"CC",x"CC",x"CC",x"7C",x"00",x"00",x"00",x"78",x"CC",x"FC",x"C0",x"78",x"00",x"00",x"00",x"78",x"CC",x"FC",x"C0",x"78",x"00",x"1C",x"30",x"30",x"78",x"30",x"30",x"30",x"00",x"1C",x"30",x"30",x"78",x"30",x"30",x"30",x"00",x"00",x"00",x"7C",x"CC",x"CC",x"7C",x"0C",x"78",x"00",x"00",x"7C",x"CC",x"CC",x"7C",x"0C",x"78",
															x"C0",x"C0",x"F8",x"CC",x"CC",x"CC",x"CC",x"00",x"C0",x"C0",x"F8",x"CC",x"CC",x"CC",x"CC",x"00",x"00",x"30",x"00",x"30",x"30",x"30",x"30",x"00",x"00",x"30",x"00",x"30",x"30",x"30",x"30",x"00",x"00",x"18",x"00",x"18",x"18",x"18",x"18",x"70",x"00",x"18",x"00",x"18",x"18",x"18",x"18",x"70",x"C0",x"C0",x"CC",x"D8",x"F0",x"D8",x"CC",x"00",x"C0",x"C0",x"CC",x"D8",x"F0",x"D8",x"CC",x"00",
															x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"00",x"00",x"EC",x"FE",x"D6",x"D6",x"D6",x"00",x"00",x"00",x"EC",x"FE",x"D6",x"D6",x"D6",x"00",x"00",x"00",x"D8",x"EC",x"CC",x"CC",x"CC",x"00",x"00",x"00",x"D8",x"EC",x"CC",x"CC",x"CC",x"00",x"00",x"00",x"3C",x"66",x"66",x"66",x"3C",x"00",x"00",x"00",x"3C",x"66",x"66",x"66",x"3C",x"00",
															x"00",x"00",x"F8",x"CC",x"CC",x"F8",x"C0",x"C0",x"00",x"00",x"F8",x"CC",x"CC",x"F8",x"C0",x"C0",x"00",x"00",x"7C",x"CC",x"CC",x"7C",x"0C",x"0C",x"00",x"00",x"7C",x"CC",x"CC",x"7C",x"0C",x"0C",x"00",x"00",x"D8",x"EC",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"D8",x"EC",x"C0",x"C0",x"C0",x"00",x"00",x"00",x"78",x"C0",x"78",x"0C",x"F8",x"00",x"00",x"00",x"78",x"C0",x"78",x"0C",x"F8",x"00",
															x"00",x"30",x"7C",x"30",x"30",x"30",x"1C",x"00",x"00",x"30",x"7C",x"30",x"30",x"30",x"1C",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"DC",x"6C",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"DC",x"6C",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"78",x"30",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"78",x"30",x"00",x"00",x"00",x"D6",x"D6",x"D6",x"FE",x"6C",x"00",x"00",x"00",x"D6",x"D6",x"D6",x"FE",x"6C",x"00",
															x"00",x"00",x"CC",x"78",x"30",x"78",x"CC",x"00",x"00",x"00",x"CC",x"78",x"30",x"78",x"CC",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"7C",x"0C",x"78",x"00",x"00",x"CC",x"CC",x"CC",x"7C",x"0C",x"78",x"00",x"00",x"FC",x"18",x"30",x"60",x"FC",x"00",x"00",x"00",x"FC",x"18",x"30",x"60",x"FC",x"00",x"0E",x"18",x"18",x"30",x"18",x"18",x"0E",x"00",x"0E",x"18",x"18",x"30",x"18",x"18",x"0E",x"00",
															x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"70",x"18",x"18",x"0C",x"18",x"18",x"70",x"00",x"70",x"18",x"18",x"0C",x"18",x"18",x"70",x"00",x"60",x"F2",x"9E",x"0C",x"00",x"00",x"00",x"00",x"60",x"F2",x"9E",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
															x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF");												
	
	constant HYDLIDE_CHR_ROM : CHR_ROM_ARRAY := (x"08", x"2C", x"29", x"23", x"26", x"26", x"23", x"21", x"09", x"0F", x"0F", x"06", x"05", x"05", x"00", x"12", x"C4", x"CC", x"64", x"F0", x"D8", x"D8", x"F8", x"E0", x"64", x"7C", x"FC", x"18", x"28", x"28", x"08", x"1E", x"72", x"01", x"00", x"00", x"00", x"07", x"07", x"00", x"77", x"3F", x"37", x"07", x"07", x"07", x"07", x"00", x"9C", x"B6", x"A2", x"B6", x"5C", x"60", x"70", x"70", x"E2", x"DD", x"DD", x"DD", x"E2", x"7C", x"70", x"70", x"03", x"8B", x"84", x"4E", x"4B", x"2B", x"2E", x"04", x"04", x"07", x"0F", x"03", x"05", x"05", x"11", x"13", x"A0", x"60", x"60", x"80", x"80", x"90", x"E0", x"00", x"20", x"E0", x"E0", x"F0", x"F0", x"F0", x"E0", x"E0", x"05", x"28", x"2C", x"24", x"68", x"68", x"3C", x"1C", x"17", x"17", x"17", x"17", x"5F", x"7E", x"3C", x"1C", x"E0", x"00", x"00", x"00", x"10", x"18", x"38", x"70", x"E0", x"E0", x"E0", x"E0", x"F0", x"78", x"38", x"70", 
															x"08", x"0D", x"0E", x"00", x"04", x"04", x"02", x"01", x"09", x"0E", x"0D", x"07", x"07", x"07", x"03", x"1B", x"C4", x"CE", x"CE", x"C2", x"CA", x"CA", x"12", x"E2", x"44", x"7C", x"7C", x"78", x"78", x"78", x"F0", x"E0", x"1A", x"21", x"20", x"38", x"18", x"07", x"07", x"00", x"27", x"5F", x"5F", x"5F", x"27", x"1F", x"07", x"00", x"17", x"E0", x"00", x"00", x"70", x"70", x"70", x"70", x"F7", x"FE", x"F6", x"F0", x"F0", x"70", x"70", x"70", x"11", x"19", x"12", x"47", x"4D", x"4D", x"47", x"43", x"12", x"1E", x"1F", x"0C", x"0A", x"0A", x"00", x"04", x"88", x"98", x"C8", x"E0", x"B0", x"B0", x"C0", x"B8", x"C8", x"F8", x"F8", x"30", x"50", x"50", x"3C", x"46", x"45", x"43", x"E1", x"01", x"0E", x"0E", x"0E", x"0E", x"0F", x"0F", x"FF", x"6F", x"6F", x"0E", x"0E", x"0E", x"6C", x"44", x"6C", x"38", x"C0", x"E0", x"E0", x"00", x"BA", x"BA", x"BA", x"C4", x"F8", x"E0", x"E0", x"00", 
															x"03", x"0B", x"04", x"8E", x"8B", x"4B", x"6E", x"24", x"04", x"07", x"0F", x"03", x"05", x"15", x"11", x"13", x"A0", x"60", x"60", x"80", x"80", x"90", x"E0", x"00", x"20", x"E0", x"E0", x"F0", x"F0", x"F0", x"E0", x"E0", x"25", x"28", x"2C", x"24", x"00", x"00", x"03", x"07", x"17", x"17", x"17", x"17", x"13", x"01", x"03", x"07", x"E0", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"11", x"1B", x"1D", x"01", x"09", x"09", x"04", x"33", x"12", x"1C", x"1A", x"0E", x"0E", x"0E", x"37", x"47", x"88", x"98", x"98", x"84", x"94", x"94", x"24", x"C4", x"88", x"F8", x"F8", x"E0", x"F0", x"F0", x"E0", x"C0", x"44", x"43", x"70", x"30", x"0E", x"0E", x"0E", x"0E", x"BF", x"BF", x"BF", x"4F", x"3F", x"0E", x"0E", x"0E", x"44", x"84", x"0E", x"00", x"00", x"E0", x"E0", x"00", x"E0", x"E0", x"EE", x"FC", x"EC", x"E0", x"E0", x"00", 
															x"05", x"29", x"21", x"27", x"21", x"31", x"39", x"7C", x"07", x"2F", x"2F", x"28", x"2F", x"2F", x"27", x"0B", x"00", x"00", x"00", x"C0", x"00", x"18", x"38", x"70", x"C0", x"E0", x"E0", x"20", x"E0", x"E0", x"C0", x"A0", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"64", x"65", x"0C", x"06", x"02", x"1C", x"1C", x"00", x"EF", x"E9", x"E9", x"E9", x"86", x"00", x"00", x"00", x"50", x"56", x"66", x"C6", x"F0", x"70", x"70", x"70", x"04", x"88", x"88", x"4F", x"48", x"28", x"38", x"71", x"07", x"8F", x"8F", x"48", x"4F", x"2F", x"2F", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"F0", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"80", x"00", x"33", x"13", x"13", x"13", x"13", x"01", x"00", x"00", x"00", x"2C", x"2F", x"20", x"03", x"1E", x"0E", x"06", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"60", x"80", x"E0", x"20", x"C0", x"18", x"38", x"70", 
															x"04", x"08", x"00", x"00", x"00", x"30", x"3F", x"1F", x"07", x"0F", x"0F", x"0F", x"0F", x"0F", x"03", x"2D", x"00", x"02", x"02", x"02", x"02", x"1A", x"FA", x"FF", x"C0", x"E2", x"E2", x"E2", x"E2", x"E2", x"82", x"60", x"1F", x"7F", x"6F", x"7F", x"0F", x"00", x"00", x"00", x"F1", x"81", x"8F", x"83", x"61", x"1C", x"1C", x"00", x"F0", x"E0", x"E0", x"E0", x"80", x"00", x"00", x"00", x"16", x"06", x"E0", x"80", x"70", x"70", x"70", x"70", x"0F", x"0F", x"0F", x"0F", x"03", x"00", x"00", x"00", x"65", x"65", x"0C", x"06", x"1E", x"1C", x"1C", x"1C", x"E0", x"EF", x"E9", x"E9", x"E9", x"06", x"00", x"00", x"40", x"50", x"76", x"D6", x"86", x"70", x"70", x"00", x"03", x"33", x"13", x"13", x"13", x"11", x"00", x"00", x"00", x"00", x"2F", x"2C", x"23", x"02", x"01", x"03", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"60", x"80", x"E0", x"20", x"C0", x"00", x"C0", x"C0", 
															x"1F", x"1F", x"6F", x"6F", x"63", x"00", x"00", x"00", x"11", x"E1", x"8F", x"83", x"9D", x"7C", x"1C", x"1C", x"F0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"16", x"06", x"E0", x"80", x"00", x"70", x"70", x"00", x"03", x"05", x"05", x"02", x"0C", x"1B", x"0F", x"16", x"03", x"06", x"06", x"01", x"09", x"16", x"10", x"25", x"80", x"40", x"40", x"80", x"A0", x"D0", x"B0", x"D8", x"00", x"80", x"80", x"00", x"30", x"28", x"48", x"00", x"33", x"63", x"42", x"03", x"13", x"01", x"02", x"07", x"2A", x"4A", x"21", x"52", x"42", x"02", x"43", x"06", x"58", x"CC", x"AC", x"C0", x"20", x"68", x"30", x"00", x"90", x"28", x"40", x"A4", x"40", x"10", x"20", x"00", x"03", x"05", x"05", x"03", x"01", x"02", x"07", x"16", x"03", x"06", x"06", x"02", x"00", x"07", x"04", x"09", x"80", x"C0", x"C0", x"80", x"80", x"C0", x"80", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", 
															x"7B", x"43", x"45", x"02", x"06", x"0C", x"44", x"1C", x"20", x"5A", x"16", x"45", x"44", x"0A", x"08", x"18", x"C0", x"40", x"80", x"C0", x"60", x"60", x"30", x"40", x"00", x"80", x"40", x"A0", x"00", x"10", x"20", x"60", x"02", x"07", x"06", x"03", x"0D", x"0B", x"1E", x"17", x"03", x"04", x"05", x"02", x"09", x"16", x"11", x"24", x"80", x"C0", x"80", x"00", x"B0", x"D0", x"F0", x"98", x"00", x"00", x"40", x"80", x"20", x"28", x"08", x"40", x"33", x"63", x"43", x"03", x"03", x"01", x"02", x"07", x"0A", x"4A", x"28", x"2A", x"42", x"42", x"03", x"06", x"D8", x"4C", x"8C", x"C0", x"60", x"28", x"30", x"00", x"10", x"80", x"48", x"A4", x"40", x"50", x"20", x"00", x"13", x"17", x"06", x"02", x"1E", x"04", x"04", x"00", x"0A", x"16", x"15", x"04", x"14", x"0A", x"00", x"00", x"5C", x"CE", x"86", x"C0", x"88", x"C0", x"C0", x"40", x"90", x"14", x"45", x"8A", x"C1", x"01", x"88", x"E0", 
															x"33", x"22", x"21", x"21", x"01", x"11", x"03", x"07", x"0A", x"11", x"30", x"11", x"10", x"01", x"01", x"00", x"C0", x"C0", x"00", x"80", x"80", x"00", x"80", x"80", x"00", x"00", x"80", x"00", x"00", x"80", x"00", x"00", x"13", x"13", x"03", x"06", x"1E", x"0A", x"04", x"00", x"0A", x"12", x"14", x"04", x"14", x"04", x"00", x"00", x"DC", x"4E", x"82", x"C0", x"80", x"C0", x"C0", x"40", x"10", x"94", x"5D", x"92", x"C2", x"10", x"82", x"E0", x"07", x"0F", x"13", x"15", x"35", x"35", x"39", x"3E", x"00", x"00", x"0C", x"0E", x"0E", x"0E", x"06", x"01", x"E0", x"F0", x"C8", x"A8", x"AC", x"AC", x"9C", x"7C", x"00", x"00", x"30", x"70", x"70", x"70", x"60", x"80", x"5D", x"5E", x"5F", x"B7", x"9D", x"7B", x"0C", x"00", x"03", x"01", x"40", x"00", x"00", x"31", x"00", x"00", x"BC", x"7C", x"FA", x"F9", x"F6", x"B1", x"DA", x"64", x"C0", x"80", x"02", x"10", x"04", x"20", x"92", x"00", 
															x"07", x"0F", x"19", x"15", x"35", x"35", x"33", x"0F", x"00", x"00", x"06", x"0E", x"0E", x"0E", x"0C", x"30", x"E0", x"F0", x"F8", x"F8", x"FC", x"FC", x"FC", x"FC", x"00", x"C0", x"70", x"30", x"28", x"58", x"38", x"18", x"BF", x"BF", x"5B", x"A7", x"9D", x"7B", x"0C", x"00", x"38", x"00", x"41", x"03", x"0C", x"31", x"00", x"00", x"FC", x"FC", x"FA", x"D9", x"F6", x"B1", x"DA", x"66", x"38", x"70", x"F2", x"C0", x"04", x"20", x"12", x"00", x"07", x"0F", x"1B", x"17", x"37", x"3F", x"3F", x"3F", x"00", x"00", x"04", x"08", x"08", x"00", x"01", x"04", x"E0", x"F0", x"F8", x"F8", x"FC", x"FC", x"FC", x"FC", x"00", x"C0", x"E0", x"70", x"B0", x"38", x"78", x"28", x"5F", x"5F", x"5F", x"B7", x"9D", x"7B", x"0C", x"00", x"00", x"04", x"4D", x"03", x"0C", x"31", x"00", x"00", x"FC", x"FC", x"7A", x"D9", x"F6", x"B1", x"DA", x"64", x"F8", x"F8", x"72", x"C0", x"04", x"20", x"12", x"00", 
															x"3B", x"37", x"58", x"9B", x"6F", x"8D", x"5B", x"26", x"07", x"0F", x"47", x"03", x"20", x"04", x"48", x"00", x"DA", x"EA", x"1A", x"ED", x"B9", x"DE", x"30", x"00", x"E0", x"F0", x"F2", x"C0", x"30", x"8C", x"00", x"00", x"37", x"3B", x"03", x"9B", x"6F", x"8D", x"5B", x"26", x"38", x"3C", x"3C", x"00", x"20", x"04", x"48", x"00", x"F9", x"FA", x"FA", x"ED", x"B9", x"DE", x"30", x"00", x"30", x"70", x"B2", x"C0", x"30", x"8C", x"00", x"00", x"3F", x"3F", x"5F", x"9F", x"6F", x"8D", x"5B", x"26", x"00", x"00", x"44", x"0D", x"23", x"04", x"48", x"00", x"FA", x"FA", x"7A", x"ED", x"B9", x"DE", x"30", x"00", x"E8", x"F0", x"62", x"48", x"30", x"8C", x"00", x"00", x"03", x"27", x"29", x"29", x"2B", x"2F", x"25", x"00", x"00", x"20", x"26", x"26", x"24", x"20", x"22", x"73", x"80", x"C0", x"20", x"20", x"A0", x"E0", x"40", x"00", x"80", x"40", x"E0", x"E0", x"60", x"20", x"C0", x"80", 
															x"37", x"31", x"07", x"05", x"03", x"0E", x"0A", x"00", x"10", x"12", x"00", x"02", x"00", x"02", x"06", x"00", x"DE", x"12", x"D2", x"52", x"EC", x"E0", x"E0", x"A0", x"C0", x"8C", x"CC", x"CC", x"00", x"00", x"00", x"60", x"07", x"4F", x"49", x"29", x"2D", x"1F", x"1A", x"00", x"00", x"40", x"46", x"26", x"22", x"10", x"15", x"39", x"00", x"40", x"A0", x"A0", x"E0", x"00", x"C0", x"80", x"80", x"80", x"40", x"40", x"00", x"C0", x"00", x"40", x"0B", x"08", x"0B", x"0A", x"09", x"1C", x"14", x"0C", x"10", x"11", x"10", x"11", x"00", x"00", x"08", x"00", x"C0", x"80", x"E0", x"A0", x"C4", x"0C", x"14", x"18", x"00", x"40", x"00", x"40", x"00", x"00", x"08", x"00", x"02", x"05", x"0D", x"0E", x"0E", x"0F", x"03", x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"03", x"80", x"C8", x"E8", x"E8", x"E8", x"E8", x"88", x"00", x"80", x"48", x"28", x"28", x"28", x"28", x"88", x"9C", 
															x"F7", x"D9", x"D7", x"F5", x"63", x"0E", x"0A", x"00", x"F0", x"A2", x"A0", x"92", x"60", x"02", x"06", x"00", x"D8", x"18", x"C0", x"40", x"E0", x"E0", x"E0", x"A0", x"C8", x"88", x"C0", x"C0", x"00", x"00", x"00", x"60", x"37", x"31", x"07", x"05", x"0F", x"0E", x"0E", x"0A", x"10", x"12", x"00", x"02", x"00", x"00", x"00", x"06", x"C0", x"1E", x"D2", x"52", x"92", x"EC", x"A0", x"00", x"C0", x"80", x"CC", x"CC", x"8C", x"00", x"60", x"00", x"03", x"08", x"0B", x"0A", x"09", x"08", x"01", x"03", x"00", x"11", x"10", x"11", x"10", x"00", x"00", x"00", x"C0", x"80", x"E0", x"A0", x"C0", x"00", x"C0", x"40", x"00", x"40", x"00", x"40", x"00", x"00", x"00", x"80", x"07", x"F9", x"D7", x"D5", x"FF", x"6E", x"0E", x"0A", x"00", x"F2", x"A0", x"A2", x"90", x"60", x"00", x"06", x"D8", x"18", x"C0", x"40", x"80", x"E0", x"A0", x"00", x"C8", x"88", x"C0", x"C0", x"80", x"00", x"60", x"00", 
															x"08", x"0E", x"0F", x"E9", x"62", x"20", x"23", x"34", x"00", x"00", x"00", x"F6", x"EF", x"E7", x"45", x"47", x"10", x"70", x"F0", x"90", x"40", x"00", x"C0", x"38", x"00", x"00", x"00", x"68", x"F0", x"E0", x"A0", x"F0", x"3E", x"1F", x"3F", x"FF", x"7F", x"39", x"19", x"00", x"03", x"01", x"30", x"F9", x"7C", x"3F", x"1F", x"00", x"78", x"FC", x"E4", x"E0", x"F8", x"FC", x"FE", x"00", x"C0", x"80", x"18", x"98", x"38", x"9C", x"8E", x"70", x"00", x"01", x"07", x"7C", x"72", x"30", x"16", x"30", x"00", x"00", x"00", x"73", x"7F", x"7F", x"65", x"07", x"40", x"E0", x"E0", x"E8", x"48", x"38", x"70", x"E0", x"00", x"00", x"00", x"08", x"A8", x"D8", x"B0", x"80", x"39", x"1F", x"03", x"03", x"03", x"0E", x"04", x"00", x"07", x"00", x"00", x"03", x"00", x"10", x"18", x"0C", x"F0", x"FF", x"FE", x"FE", x"FC", x"3C", x"08", x"00", x"F0", x"FF", x"7E", x"BE", x"1C", x"02", x"06", x"0C", 
															x"08", x"0E", x"0F", x"0F", x"03", x"00", x"00", x"07", x"00", x"00", x"00", x"10", x"0C", x"07", x"03", x"04", x"10", x"70", x"F0", x"F7", x"C6", x"04", x"0C", x"FE", x"00", x"00", x"00", x"0F", x"37", x"E7", x"C2", x"18", x"07", x"0F", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"06", x"0F", x"0F", x"1F", x"1F", x"3F", x"3F", x"0E", x"FC", x"F8", x"FC", x"FE", x"FF", x"CE", x"C8", x"00", x"78", x"F8", x"FC", x"FE", x"FF", x"FE", x"F8", x"00", x"3E", x"1F", x"0F", x"1F", x"1F", x"3F", x"7F", x"00", x"03", x"01", x"00", x"19", x"1C", x"39", x"71", x"0E", x"78", x"FC", x"FF", x"F9", x"FC", x"9C", x"90", x"00", x"C0", x"80", x"13", x"9F", x"3E", x"FC", x"F0", x"00", x"39", x"1F", x"03", x"03", x"03", x"01", x"00", x"00", x"07", x"01", x"00", x"03", x"00", x"00", x"01", x"03", x"E0", x"E0", x"E0", x"F0", x"F8", x"F8", x"BC", x"00", x"E0", x"E0", x"E0", x"F0", x"78", x"78", x"3C", x"80", 
															x"0F", x"1F", x"3F", x"FF", x"7F", x"33", x"03", x"00", x"0E", x"1F", x"3F", x"FF", x"7F", x"3F", x"0F", x"00", x"FC", x"F8", x"F8", x"FC", x"FC", x"FC", x"FC", x"00", x"78", x"F8", x"F8", x"FC", x"FC", x"FC", x"FC", x"38", x"00", x"0F", x"18", x"30", x"20", x"02", x"8F", x"78", x"0F", x"30", x"67", x"4F", x"DF", x"FF", x"FF", x"78", x"00", x"80", x"20", x"10", x"0C", x"60", x"F0", x"1C", x"00", x"00", x"C0", x"E0", x"F0", x"FE", x"FE", x"1C", x"04", x"3C", x"14", x"3C", x"19", x"5E", x"1E", x"3A", x"40", x"40", x"40", x"40", x"21", x"22", x"E4", x"88", x"04", x"0C", x"8E", x"9E", x"9C", x"4C", x"5E", x"5E", x"00", x"10", x"A0", x"A0", x"80", x"50", x"60", x"60", x"02", x"0E", x"1E", x"9E", x"4C", x"0E", x"0F", x"0D", x"20", x"30", x"20", x"A0", x"50", x"30", x"70", x"50", x"07", x"08", x"12", x"0B", x"27", x"17", x"1F", x"15", x"00", x"07", x"08", x"10", x"10", x"20", x"20", x"20", 
															x"80", x"60", x"10", x"90", x"A0", x"F0", x"D0", x"50", x"00", x"80", x"E0", x"20", x"10", x"08", x"08", x"08", x"35", x"1F", x"1D", x"1F", x"1D", x"0F", x"1B", x"0F", x"00", x"0F", x"05", x"07", x"05", x"07", x"83", x"27", x"78", x"F8", x"D8", x"F8", x"D0", x"F8", x"B0", x"E0", x"00", x"E0", x"C0", x"E0", x"C0", x"C0", x"82", x"C8", x"00", x"00", x"42", x"42", x"24", x"00", x"54", x"00", x"3C", x"7E", x"FF", x"FF", x"FF", x"FF", x"2A", x"7E", x"3C", x"00", x"3C", x"00", x"BC", x"01", x"3C", x"82", x"42", x"7E", x"42", x"7E", x"42", x"7E", x"00", x"00", x"00", x"08", x"08", x"10", x"00", x"A8", x"00", x"10", x"3C", x"7E", x"FE", x"FF", x"FF", x"57", x"7F", x"0F", x"00", x"18", x"00", x"18", x"00", x"18", x"40", x"11", x"1F", x"07", x"1F", x"07", x"1F", x"07", x"0E", x"00", x"00", x"20", x"40", x"40", x"00", x"00", x"20", x"20", x"3C", x"5E", x"BF", x"BF", x"FF", x"FF", x"5E", x"5E", 
															x"20", x"20", x"20", x"20", x"80", x"21", x"00", x"8A", x"5E", x"5E", x"5E", x"5E", x"7E", x"5E", x"3C", x"00", x"00", x"00", x"31", x"7B", x"4F", x"0F", x"1B", x"13", x"01", x"03", x"37", x"7F", x"4D", x"0D", x"1F", x"1F", x"00", x"00", x"80", x"C0", x"E0", x"E0", x"C0", x"C0", x"80", x"C0", x"E0", x"F0", x"B8", x"B8", x"FC", x"FC", x"1D", x"1C", x"18", x"10", x"10", x"10", x"17", x"00", x"27", x"27", x"2F", x"3F", x"1F", x"1F", x"17", x"00", x"B8", x"38", x"1C", x"0C", x"04", x"70", x"70", x"70", x"CE", x"CE", x"FE", x"FE", x"FE", x"FC", x"70", x"70", x"00", x"00", x"70", x"C6", x"9F", x"9E", x"5E", x"1C", x"01", x"07", x"7F", x"DF", x"97", x"97", x"5F", x"1F", x"00", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"20", x"3C", x"3C", x"06", x"63", x"78", x"3C", x"18", x"2F", x"27", x"27", x"1F", x"7F", x"7F", x"3C", x"18", 
															x"00", x"00", x"00", x"00", x"28", x"CC", x"3C", x"38", x"F0", x"F8", x"F8", x"F8", x"F8", x"FC", x"FC", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"CC", x"3E", x"02", x"00", x"08", x"08", x"80", x"C0", x"EC", x"FE", x"F2", x"F0", x"F8", x"F8", x"08", x"10", x"10", x"10", x"20", x"0E", x"0E", x"0E", x"7F", x"7F", x"7F", x"7F", x"3F", x"0F", x"0E", x"0E", x"00", x"00", x"20", x"20", x"20", x"08", x"E8", x"00", x"F8", x"FC", x"FC", x"FC", x"FC", x"F8", x"E8", x"00", x"1D", x"1C", x"18", x"10", x"10", x"17", x"17", x"07", x"27", x"27", x"2F", x"3F", x"1F", x"1F", x"17", x"07", x"80", x"38", x"3C", x"0C", x"0C", x"04", x"70", x"00", x"FE", x"CE", x"CE", x"FE", x"FE", x"FE", x"7C", x"00", x"18", x"1C", x"3C", x"26", x"23", x"20", x"03", x"07", x"1F", x"07", x"27", x"2F", x"2F", x"2F", x"0F", x"07", 
															x"00", x"00", x"00", x"00", x"20", x"C0", x"80", x"C0", x"F0", x"F0", x"F0", x"F8", x"F8", x"FC", x"FC", x"C0", x"04", x"04", x"08", x"08", x"10", x"00", x"0E", x"00", x"3F", x"7F", x"7F", x"7F", x"3F", x"0F", x"0E", x"00", x"00", x"00", x"10", x"10", x"10", x"E0", x"E8", x"E0", x"F8", x"FC", x"FC", x"FC", x"FC", x"F8", x"E8", x"E0", x"00", x"00", x"03", x"05", x"0D", x"33", x"37", x"B7", x"00", x"1F", x"3C", x"7A", x"72", x"4C", x"48", x"48", x"00", x"20", x"38", x"7C", x"7E", x"FE", x"FE", x"FE", x"80", x"C0", x"D8", x"A8", x"AA", x"1A", x"1A", x"1E", x"56", x"66", x"66", x"66", x"E6", x"E6", x"1C", x"01", x"A9", x"99", x"99", x"B9", x"7B", x"BF", x"0F", x"01", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"FF", x"FE", x"33", x"2B", x"2B", x"89", x"89", x"8B", x"2F", x"FE", x"17", x"2A", x"1D", x"3F", x"3B", x"53", x"3F", x"5F", x"17", x"2A", x"1D", x"3F", x"3B", x"53", x"36", x"58", 
															x"E4", x"FA", x"FC", x"FE", x"FC", x"FE", x"FC", x"FE", x"E4", x"C2", x"E0", x"68", x"A0", x"C8", x"54", x"28", x"2E", x"37", x"1B", x"0E", x"02", x"06", x"1C", x"0F", x"2C", x"1E", x"04", x"01", x"01", x"07", x"1B", x"08", x"FE", x"EE", x"DC", x"FC", x"30", x"3C", x"1E", x"FE", x"40", x"D4", x"E0", x"04", x"D0", x"C4", x"E0", x"02", x"1E", x"7C", x"F8", x"FD", x"FB", x"C1", x"81", x"01", x"02", x"00", x"00", x"00", x"00", x"03", x"03", x"01", x"78", x"3E", x"1F", x"BF", x"DF", x"83", x"81", x"80", x"40", x"00", x"00", x"00", x"00", x"C0", x"C0", x"80", x"18", x"38", x"7D", x"7F", x"7D", x"71", x"61", x"20", x"08", x"00", x"00", x"00", x"03", x"03", x"01", x"00", x"18", x"1C", x"BE", x"FE", x"BE", x"8E", x"86", x"04", x"10", x"00", x"00", x"00", x"C0", x"C0", x"80", x"00", x"C3", x"E7", x"66", x"A5", x"5A", x"00", x"3C", x"00", x"C3", x"E7", x"66", x"BD", x"42", x"24", x"00", x"18", 
															x"00", x"24", x"5A", x"C3", x"BD", x"42", x"81", x"00", x"00", x"3C", x"42", x"E7", x"81", x"5A", x"81", x"00", x"00", x"00", x"04", x"02", x"06", x"0D", x"16", x"11", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"07", x"00", x"00", x"C0", x"20", x"20", x"30", x"54", x"94", x"00", x"00", x"00", x"00", x"40", x"C0", x"E0", x"E0", x"0B", x"0C", x"15", x"12", x"09", x"00", x"00", x"00", x"07", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"C8", x"90", x"70", x"68", x"30", x"80", x"00", x"00", x"F0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"06", x"01", x"1F", x"25", x"08", x"15", x"33", x"00", x"00", x"00", x"00", x"03", x"07", x"0B", x"0F", x"00", x"C0", x"68", x"A4", x"B4", x"DC", x"0C", x"B8", x"00", x"00", x"00", x"00", x"40", x"A0", x"F0", x"E0", x"29", x"46", x"18", x"19", x"0E", x"0B", x"09", x"04", x"07", x"0B", x"07", x"07", x"01", x"00", x"00", x"00", 
															x"A2", x"5C", x"98", x"74", x"F8", x"80", x"E0", x"00", x"D0", x"E0", x"60", x"80", x"00", x"00", x"00", x"00", x"10", x"08", x"18", x"7D", x"BE", x"18", x"10", x"08", x"10", x"08", x"18", x"65", x"AE", x"18", x"10", x"08", x"04", x"32", x"9A", x"3C", x"79", x"8D", x"40", x"24", x"04", x"32", x"8A", x"24", x"59", x"8D", x"40", x"24", x"00", x"01", x"3E", x"00", x"17", x"02", x"19", x"0D", x"0C", x"11", x"0F", x"03", x"14", x"7D", x"E6", x"CE", x"00", x"3F", x"FF", x"3F", x"FF", x"1E", x"00", x"00", x"3F", x"C0", x"00", x"C0", x"E3", x"31", x"7F", x"FF", x"00", x"C0", x"E0", x"F0", x"FA", x"C1", x"01", x"01", x"E0", x"38", x"E0", x"00", x"30", x"C0", x"F2", x"FE", x"0C", x"1C", x"76", x"03", x"00", x"00", x"00", x"14", x"03", x"03", x"01", x"00", x"07", x"0F", x"1C", x"28", x"00", x"26", x"C7", x"9F", x"BE", x"80", x"08", x"00", x"FF", x"F9", x"78", x"E4", x"C9", x"F0", x"30", x"00", 
															x"72", x"2C", x"00", x"00", x"88", x"00", x"04", x"00", x"CC", x"E0", x"E0", x"F8", x"F0", x"18", x"08", x"00", x"00", x"00", x"00", x"00", x"14", x"01", x"18", x"0C", x"00", x"00", x"03", x"00", x"14", x"3D", x"66", x"FE", x"00", x"00", x"00", x"00", x"0F", x"07", x"00", x"00", x"00", x"00", x"FF", x"FF", x"3F", x"38", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"E1", x"00", x"01", x"00", x"00", x"00", x"F0", x"F8", x"E0", x"E1", x"F2", x"7C", x"7C", x"06", x"03", x"00", x"00", x"00", x"05", x"F3", x"03", x"01", x"00", x"03", x"03", x"07", x"02", x"00", x"26", x"C7", x"9F", x"BE", x"80", x"40", x"00", x"FF", x"F9", x"78", x"E4", x"C9", x"F0", x"30", x"00", x"61", x"32", x"0C", x"80", x"80", x"00", x"10", x"00", x"DE", x"EC", x"E0", x"F8", x"F8", x"38", x"20", x"00", x"00", x"08", x"18", x"38", x"39", x"79", x"7B", x"7B", x"00", x"08", x"00", x"00", x"00", x"00", x"04", x"04", 
															x"80", x"C1", x"41", x"63", x"77", x"B6", x"B6", x"B6", x"00", x"00", x"00", x"00", x"88", x"6B", x"7F", x"5D", x"80", x"98", x"0C", x"0E", x"1E", x"3E", x"9F", x"EF", x"00", x"10", x"00", x"00", x"00", x"00", x"60", x"10", x"F7", x"EE", x"D0", x"D5", x"D5", x"E8", x"F8", x"F8", x"08", x"11", x"2F", x"3F", x"3F", x"1E", x"04", x"04", x"B6", x"D5", x"DD", x"EB", x"76", x"7E", x"BC", x"98", x"49", x"2A", x"22", x"14", x"89", x"81", x"43", x"67", x"F7", x"7B", x"19", x"5D", x"5C", x"5F", x"37", x"25", x"08", x"84", x"E6", x"A2", x"A3", x"AD", x"FD", x"FF", x"7C", x"7C", x"75", x"31", x"31", x"31", x"12", x"02", x"00", x"00", x"08", x"08", x"08", x"09", x"0A", x"0A", x"C1", x"C3", x"87", x"C1", x"C1", x"E1", x"A1", x"80", x"3E", x"04", x"40", x"02", x"03", x"21", x"A1", x"80", x"0F", x"9F", x"97", x"C6", x"D6", x"D6", x"04", x"00", x"30", x"20", x"28", x"78", x"58", x"58", x"08", x"08", 
															x"00", x"01", x"03", x"07", x"07", x"0E", x"0D", x"1B", x"00", x"01", x"00", x"00", x"00", x"01", x"02", x"04", x"80", x"C1", x"41", x"63", x"77", x"14", x"00", x"22", x"00", x"00", x"80", x"80", x"88", x"EB", x"FF", x"DD", x"80", x"E0", x"30", x"38", x"38", x"9C", x"EC", x"E4", x"00", x"40", x"80", x"80", x"80", x"60", x"10", x"18", x"1B", x"1B", x"1B", x"16", x"17", x"0F", x"15", x"15", x"04", x"04", x"04", x"09", x"08", x"14", x"1F", x"1F", x"B6", x"D5", x"5D", x"6B", x"76", x"7E", x"BC", x"98", x"49", x"2A", x"A2", x"94", x"89", x"81", x"43", x"67", x"F6", x"7A", x"1A", x"7E", x"5E", x"1E", x"1E", x"3E", x"08", x"84", x"FE", x"EA", x"EA", x"E0", x"E0", x"C0", x"0E", x"0C", x"0B", x"0B", x"05", x"05", x"00", x"00", x"01", x"03", x"04", x"04", x"07", x"07", x"00", x"00", x"C3", x"E3", x"C1", x"C1", x"41", x"41", x"01", x"01", x"3C", x"00", x"00", x"40", x"C0", x"C1", x"01", x"01", 
															x"BE", x"BE", x"96", x"C4", x"C4", x"E8", x"F0", x"50", x"40", x"40", x"68", x"28", x"28", x"40", x"50", x"70", x"08", x"0F", x"0E", x"07", x"0A", x"07", x"08", x"1F", x"04", x"00", x"07", x"08", x"05", x"00", x"07", x"04", x"20", x"E0", x"E0", x"C3", x"AF", x"CF", x"03", x"E0", x"40", x"00", x"C0", x"26", x"4E", x"0E", x"C6", x"24", x"2F", x"33", x"03", x"03", x"06", x"06", x"06", x"00", x"12", x"01", x"02", x"01", x"00", x"00", x"00", x"06", x"F0", x"DC", x"CC", x"C0", x"00", x"60", x"00", x"00", x"44", x"80", x"40", x"84", x"04", x"00", x"60", x"00", x"00", x"03", x"03", x"C7", x"E5", x"E7", x"60", x"03", x"00", x"00", x"07", x"60", x"62", x"60", x"33", x"12", x"40", x"C0", x"E0", x"E0", x"60", x"C0", x"00", x"C0", x"80", x"00", x"00", x"00", x"80", x"00", x"C0", x"00", x"07", x"1D", x"1B", x"03", x"13", x"18", x"0C", x"00", x"08", x"02", x"06", x"02", x"00", x"00", x"10", x"0C", 
															x"C0", x"C0", x"C0", x"C0", x"B0", x"30", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"60", x"04", x"07", x"07", x"C7", x"F7", x"F3", x"C0", x"07", x"02", x"00", x"00", x"60", x"70", x"70", x"63", x"20", x"10", x"F0", x"F0", x"F0", x"F0", x"E0", x"00", x"F8", x"20", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"0F", x"3B", x"33", x"03", x"00", x"06", x"00", x"00", x"20", x"00", x"00", x"20", x"20", x"00", x"06", x"00", x"FC", x"CC", x"C0", x"C0", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"1F", x"1B", x"23", x"33", x"00", x"06", x"00", x"00", x"02", x"01", x"12", x"01", x"00", x"00", x"06", x"00", x"F0", x"DC", x"CC", x"C0", x"60", x"60", x"60", x"00", x"44", x"80", x"40", x"84", x"04", x"00", x"00", x"60", x"07", x"05", x"0F", x"0F", x"03", x"01", x"03", x"00", x"08", x"02", x"02", x"02", x"00", x"00", x"00", x"03", 
															x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"0F", x"3B", x"33", x"03", x"06", x"06", x"06", x"00", x"20", x"00", x"00", x"20", x"20", x"00", x"00", x"06", x"F8", x"D8", x"CC", x"CC", x"00", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"00", x"04", x"89", x"1E", x"07", x"63", x"0C", x"39", x"7D", x"03", x"40", x"00", x"00", x"1C", x"03", x"06", x"07", x"00", x"80", x"0C", x"80", x"F0", x"6E", x"18", x"B7", x"00", x"00", x"00", x"00", x"00", x"D0", x"EC", x"EF", x"D3", x"38", x"01", x"64", x"08", x"00", x"60", x"06", x"3F", x"07", x"0E", x"10", x"06", x"00", x"00", x"00", x"7E", x"2C", x"10", x"CC", x"60", x"00", x"B0", x"00", x"F8", x"D0", x"A0", x"00", x"00", x"00", x"00", x"00", x"60", x"70", x"78", x"3B", x"39", x"1B", x"0D", x"0B", x"40", x"41", x"03", x"07", x"05", x"03", x"09", x"0B", 
															x"03", x"0F", x"1F", x"BE", x"5E", x"DC", x"A8", x"B0", x"02", x"84", x"C0", x"C0", x"60", x"E0", x"90", x"C0", x"1C", x"3C", x"3C", x"1E", x"02", x"02", x"01", x"00", x"07", x"21", x"01", x"03", x"03", x"02", x"00", x"00", x"0C", x"6E", x"2E", x"1C", x"80", x"C0", x"60", x"20", x"E8", x"F0", x"A0", x"D0", x"C0", x"C0", x"40", x"00", x"10", x"18", x"1B", x"19", x"0F", x"0D", x"0B", x"04", x"01", x"03", x"07", x"05", x"03", x"09", x"0B", x"07", x"08", x"18", x"B8", x"58", x"D0", x"A0", x"B0", x"08", x"80", x"C0", x"C0", x"60", x"E0", x"80", x"C0", x"E0", x"0C", x"0C", x"06", x"02", x"02", x"01", x"00", x"00", x"01", x"01", x"03", x"03", x"02", x"00", x"00", x"00", x"6C", x"2C", x"18", x"80", x"C0", x"60", x"20", x"00", x"F0", x"A0", x"D0", x"C0", x"C0", x"40", x"00", x"00", x"00", x"04", x"20", x"18", x"BE", x"0D", x"40", x"02", x"00", x"0C", x"60", x"2B", x"7E", x"15", x"40", x"06", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"80", x"3A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"02", x"00", x"07", x"8A", x"CF", x"CA", x"C7", x"C0", x"00", x"07", x"08", x"97", x"F7", x"F7", x"C8", x"C7", x"6C", x"6D", x"39", x"A1", x"96", x"A7", x"18", x"00", x"17", x"16", x"CE", x"7E", x"7E", x"7F", x"BC", x"00", x"10", x"22", x"4C", x"48", x"90", x"90", x"90", x"90", x"00", x"02", x"0C", x"09", x"11", x"12", x"12", x"12", x"00", x"00", x"00", x"10", x"20", x"24", x"48", x"48", x"00", x"00", x"80", x"80", x"00", x"04", x"09", x"0A", 
															x"90", x"90", x"90", x"90", x"48", x"4C", x"22", x"10", x"12", x"12", x"12", x"11", x"09", x"0C", x"02", x"00", x"48", x"48", x"24", x"20", x"10", x"00", x"00", x"00", x"0A", x"09", x"04", x"00", x"80", x"80", x"00", x"00", x"44", x"82", x"28", x"00", x"28", x"82", x"44", x"00", x"28", x"6C", x"C6", x"38", x"D6", x"6C", x"28", x"00", x"07", x"0F", x"1F", x"1F", x"1A", x"3A", x"3F", x"27", x"00", x"00", x"04", x"06", x"0A", x"0A", x"0F", x"17", x"00", x"80", x"C0", x"C0", x"C0", x"E0", x"E0", x"20", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"40", x"00", x"30", x"38", x"22", x"40", x"00", x"00", x"00", x"3F", x"1F", x"37", x"24", x"4F", x"1F", x"1F", x"3F", x"00", x"30", x"70", x"10", x"08", x"00", x"00", x"00", x"F0", x"E0", x"B0", x"90", x"C8", x"C0", x"E0", x"F0", x"00", x"07", x"0F", x"1F", x"1F", x"1F", x"3F", x"27", x"00", x"00", x"00", x"00", x"00", x"08", x"0E", x"17", 
															x"00", x"00", x"80", x"C0", x"C0", x"C0", x"E0", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"20", x"00", x"1C", x"0E", x"06", x"03", x"00", x"00", x"0C", x"1F", x"0F", x"0C", x"0F", x"1F", x"1F", x"3F", x"20", x"00", x"E0", x"C0", x"80", x"00", x"00", x"00", x"C0", x"E0", x"C0", x"C0", x"80", x"40", x"E0", x"F0", x"1C", x"1C", x"10", x"12", x"12", x"12", x"11", x"30", x"20", x"20", x"24", x"24", x"24", x"24", x"22", x"40", x"0E", x"0E", x"0A", x"11", x"11", x"31", x"21", x"63", x"10", x"10", x"10", x"22", x"22", x"02", x"C2", x"04", x"0C", x"0E", x"16", x"12", x"12", x"22", x"E2", x"03", x"10", x"10", x"00", x"24", x"24", x"44", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"D4", x"69", x"A0", x"C9", x"83", x"81", x"C0", x"FF", x"D4", x"69", x"A0", x"C8", x"30", x"39", x"78", x"3E", x"55", x"FA", x"F5", x"79", x"E4", x"A8", x"F2", x"74", x"04", x"5A", x"B5", x"79", x"64", x"A8", x"B2", x"74", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"04", x"40", x"00", x"02", x"00", x"08", x"00", x"FF", x"BF", x"FE", x"FF", x"EF", x"FB", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7E", x"00", x"D3", x"F7", x"F7", x"00", x"7C", x"FE", x"FE", x"AA", x"AA", x"AA", x"2A", x"0C", x"00", x"00", x"02", x"5E", x"5E", x"5E", x"DE", x"7C", x"7C", x"82", x"70", x"E8", x"E8", x"E8", x"E8", x"28", x"00", x"7C", x"8A", x"AA", x"AA", x"AA", x"AA", x"68", x"BB", x"9D", x"D4", x"B4", x"ED", x"6B", x"DE", x"BD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"40", x"02", x"10", x"00", x"00", x"08", x"FF", x"FB", x"FF", x"FF", x"FF", x"F7", x"7F", x"FF", x"FF", x"E0", x"C3", x"85", x"8D", x"B3", x"B7", x"B7", x"FF", x"FF", x"FC", x"FA", x"F2", x"CC", x"C8", x"48", x"7F", x"3F", x"27", x"57", x"55", x"E5", x"E5", x"E1", x"FF", x"DF", x"C7", x"83", x"81", x"01", x"01", x"01", x"56", x"66", x"66", x"46", x"84", x"40", x"F0", x"FE", x"A9", x"99", x"99", x"99", x"19", x"19", x"E3", x"FE", x"CC", x"D4", x"D4", x"76", x"76", x"74", x"D0", x"01", x"00", x"00", x"00", x"80", x"80", x"80", x"00", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F8", x"17", x"2A", x"1D", x"3F", x"3B", x"53", x"36", x"58", x"FF", x"C7", x"E3", x"69", x"A3", x"C9", x"57", x"29", x"E4", x"C2", x"E0", x"68", x"A0", x"C8", x"54", x"28", x"FD", x"D6", x"E0", x"F0", x"FC", x"FE", x"F8", x"F8", x"2C", x"1E", x"04", x"01", x"01", x"07", x"1B", x"08", 
															x"41", x"C5", x"C3", x"07", x"1F", x"07", x"01", x"03", x"40", x"D4", x"E0", x"04", x"D0", x"C4", x"E0", x"02", x"7F", x"80", x"BF", x"A5", x"C5", x"B9", x"A0", x"BC", x"00", x"7F", x"40", x"5B", x"3B", x"47", x"5F", x"5F", x"F8", x"00", x"F0", x"00", x"00", x"E0", x"00", x"E0", x"06", x"F3", x"0D", x"35", x"35", x"05", x"E5", x"E5", x"85", x"A1", x"A0", x"A4", x"A5", x"87", x"A0", x"40", x"43", x"5B", x"5C", x"5A", x"5B", x"5B", x"10", x"19", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"05", x"34", x"35", x"34", x"35", x"30", x"54", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7A", x"10", x"C0", x"E0", x"C0", x"20", x"00", x"00", x"A0", x"00", x"10", x"04", x"00", x"00", x"7F", x"7F", x"0E", x"18", x"0F", x"03", x"07", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"60", x"70", x"00", x"D6", x"F7", x"F7", x"00", 
															x"04", x"04", x"08", x"04", x"90", x"00", x"00", x"00", x"01", x"03", x"02", x"20", x"47", x"F3", x"B7", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E3", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E3", x"E7", x"DF", x"9F", x"1F", x"1F", x"0F", x"0F", x"0F", x"07", x"9F", x"DF", x"DF", x"5F", x"CF", x"4F", x"EE", x"64", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"68", x"F9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FD", x"4D", x"06", x"DF", x"8F", x"8F", x"27", x"27", x"61", x"20", x"A4", x"DF", x"CF", x"CF", x"C7", x"C7", x"81", x"92", x"12", x"EF", x"EF", x"E5", x"E2", x"E1", x"40", x"26", x"82", x"EE", x"C6", x"C4", x"80", x"00", x"82", x"C8", x"7C", x"2A", x"53", x"2A", x"02", x"32", x"12", x"12", x"10", x"50", x"28", x"00", x"0C", x"04", x"24", x"20", x"20", x"F8", x"78", x"1C", x"1C", x"5C", x"4C", x"54", x"48", x"07", x"07", x"01", x"02", x"83", x"83", x"83", x"83", 
															x"3C", x"28", x"14", x"01", x"35", x"29", x"15", x"09", x"C0", x"D0", x"C0", x"01", x"C1", x"D1", x"81", x"91", x"B8", x"84", x"84", x"8C", x"84", x"8C", x"84", x"8C", x"00", x"40", x"78", x"50", x"58", x"70", x"58", x"50", x"00", x"01", x"E0", x"E2", x"F2", x"F0", x"F5", x"F2", x"02", x"62", x"00", x"0C", x"0C", x"0F", x"0A", x"0D", x"05", x"C2", x"00", x"22", x"22", x"00", x"56", x"AA", x"00", x"00", x"00", x"CD", x"CC", x"FE", x"A8", x"54", x"15", x"09", x"95", x"A9", x"55", x"29", x"D5", x"69", x"E1", x"91", x"01", x"51", x"A1", x"C1", x"21", x"01", x"94", x"8D", x"95", x"8D", x"95", x"CC", x"78", x"E0", x"68", x"70", x"68", x"70", x"68", x"31", x"00", x"E0", x"F5", x"B2", x"14", x"12", x"14", x"02", x"04", x"00", x"0A", x"0D", x"6A", x"6C", x"6A", x"7C", x"0A", x"00", x"54", x"2A", x"54", x"6A", x"64", x"6A", x"64", x"00", x"A8", x"14", x"08", x"14", x"18", x"14", x"18", x"00", 
															x"14", x"10", x"0F", x"00", x"08", x"73", x"F9", x"FF", x"00", x"2E", x"10", x"00", x"27", x"04", x"02", x"FF", x"3C", x"43", x"E3", x"85", x"80", x"A6", x"82", x"00", x"3F", x"41", x"DC", x"A2", x"BE", x"80", x"BE", x"00", x"8C", x"C6", x"E3", x"67", x"FB", x"F7", x"FE", x"B9", x"F8", x"7C", x"BE", x"D8", x"46", x"59", x"46", x"39", x"AA", x"3E", x"C1", x"C9", x"C1", x"D9", x"36", x"00", x"FF", x"80", x"9C", x"C9", x"9C", x"80", x"90", x"7F", x"45", x"E1", x"45", x"65", x"73", x"41", x"C0", x"00", x"E9", x"4D", x"69", x"43", x"4D", x"72", x"4C", x"B0", x"7F", x"7F", x"7F", x"00", x"F7", x"F7", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3C", x"66", x"6E", x"76", x"66", x"66", x"3C", x"00", x"3C", x"66", x"6E", x"76", x"66", x"66", x"3C", x"00", x"08", x"18", x"38", x"18", x"18", x"18", x"18", x"00", x"08", x"18", x"38", x"18", x"18", x"18", x"18", x"00", x"3C", x"66", x"66", x"0E", x"38", x"70", x"7E", x"00", x"3C", x"66", x"66", x"0E", x"38", x"70", x"7E", x"00", x"3C", x"66", x"66", x"0C", x"66", x"66", x"3C", x"00", x"3C", x"66", x"66", x"0C", x"66", x"66", x"3C", x"00", x"0C", x"1C", x"2C", x"4C", x"7E", x"0C", x"0C", x"00", x"0C", x"1C", x"2C", x"4C", x"7E", x"0C", x"0C", x"00", x"7E", x"60", x"7C", x"06", x"66", x"66", x"3C", x"00", x"7E", x"60", x"7C", x"06", x"66", x"66", x"3C", x"00", x"3C", x"66", x"60", x"7C", x"66", x"66", x"3C", x"00", x"3C", x"66", x"60", x"7C", x"66", x"66", x"3C", x"00", x"7E", x"66", x"66", x"0C", x"18", x"18", x"18", x"00", x"7E", x"66", x"66", x"0C", x"18", x"18", x"18", x"00", 
															x"3C", x"66", x"66", x"3C", x"66", x"66", x"3C", x"00", x"3C", x"66", x"66", x"3C", x"66", x"66", x"3C", x"00", x"3C", x"66", x"66", x"3E", x"06", x"66", x"3C", x"00", x"3C", x"66", x"66", x"3E", x"06", x"66", x"3C", x"00", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"00", x"38", x"64", x"60", x"36", x"6C", x"6C", x"38", x"00", x"38", x"64", x"60", x"36", x"6C", x"6C", x"38", x"00", x"38", x"38", x"30", x"20", x"00", x"30", x"30", x"00", x"38", x"38", x"30", x"20", x"00", x"30", x"30", x"00", x"3C", x"66", x"66", x"0C", x"18", x"00", x"18", x"00", x"3C", x"66", x"66", x"0C", x"18", x"00", x"18", x"00", x"00", x"00", x"00", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"00", x"00", x"00", x"03", x"06", x"0C", x"18", x"30", x"60", x"C0", x"00", x"03", x"06", x"0C", x"18", x"30", x"60", x"C0", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"3C", x"66", x"66", x"7E", x"66", x"66", x"00", x"18", x"3C", x"66", x"66", x"7E", x"66", x"66", x"00", x"7C", x"66", x"66", x"7E", x"66", x"66", x"7C", x"00", x"7C", x"66", x"66", x"7E", x"66", x"66", x"7C", x"00", x"3C", x"66", x"60", x"60", x"60", x"66", x"3C", x"00", x"3C", x"66", x"60", x"60", x"60", x"66", x"3C", x"00", x"78", x"64", x"66", x"66", x"66", x"64", x"78", x"00", x"78", x"64", x"66", x"66", x"66", x"64", x"78", x"00", x"7E", x"60", x"60", x"7C", x"60", x"60", x"7E", x"00", x"7E", x"60", x"60", x"7C", x"60", x"60", x"7E", x"00", x"7E", x"60", x"60", x"7C", x"60", x"60", x"60", x"00", x"7E", x"60", x"60", x"7C", x"60", x"60", x"60", x"00", x"3C", x"66", x"60", x"6E", x"66", x"66", x"3C", x"00", x"3C", x"66", x"60", x"6E", x"66", x"66", x"3C", x"00", 
															x"66", x"66", x"66", x"7E", x"66", x"66", x"66", x"00", x"66", x"66", x"66", x"7E", x"66", x"66", x"66", x"00", x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"06", x"06", x"06", x"06", x"66", x"66", x"3C", x"00", x"06", x"06", x"06", x"06", x"66", x"66", x"3C", x"00", x"66", x"6C", x"78", x"70", x"78", x"6C", x"66", x"00", x"66", x"6C", x"78", x"70", x"78", x"6C", x"66", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"42", x"66", x"7E", x"66", x"66", x"66", x"66", x"00", x"42", x"66", x"7E", x"66", x"66", x"66", x"66", x"00", x"46", x"66", x"76", x"7E", x"6E", x"66", x"62", x"00", x"46", x"66", x"76", x"7E", x"6E", x"66", x"62", x"00", x"3C", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"3C", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", 
															x"7C", x"66", x"66", x"7C", x"60", x"60", x"60", x"00", x"7C", x"66", x"66", x"7C", x"60", x"60", x"60", x"00", x"3C", x"66", x"66", x"66", x"6E", x"6E", x"3E", x"00", x"3C", x"66", x"66", x"66", x"6E", x"6E", x"3E", x"00", x"7C", x"66", x"66", x"7C", x"78", x"6C", x"66", x"00", x"7C", x"66", x"66", x"7C", x"78", x"6C", x"66", x"00", x"3C", x"66", x"60", x"3C", x"06", x"66", x"3C", x"00", x"3C", x"66", x"60", x"3C", x"06", x"66", x"3C", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"66", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"66", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"66", x"66", x"66", x"66", x"66", x"3C", x"18", x"00", x"66", x"66", x"66", x"66", x"66", x"3C", x"18", x"00", x"66", x"66", x"66", x"7E", x"7E", x"66", x"42", x"00", x"66", x"66", x"66", x"7E", x"7E", x"66", x"42", x"00", 
															x"66", x"66", x"3C", x"18", x"3C", x"66", x"66", x"00", x"66", x"66", x"3C", x"18", x"3C", x"66", x"66", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"7E", x"06", x"0C", x"18", x"30", x"60", x"7E", x"00", x"7E", x"06", x"0C", x"18", x"30", x"60", x"7E", x"00", x"00", x"00", x"00", x"1F", x"1F", x"18", x"18", x"18", x"00", x"00", x"00", x"1F", x"1F", x"18", x"18", x"18", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F8", x"18", x"18", x"18", x"00", x"00", x"00", x"F8", x"F8", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"1F", x"1F", x"00", x"00", x"00", x"18", x"18", x"18", x"1F", x"1F", x"00", x"00", x"00", 
															x"18", x"18", x"18", x"F8", x"F8", x"00", x"00", x"00", x"18", x"18", x"18", x"F8", x"F8", x"00", x"00", x"00", x"18", x"3C", x"66", x"66", x"7E", x"66", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"66", x"66", x"7E", x"66", x"66", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"60", x"60", x"60", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"64", x"66", x"66", x"66", x"64", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"60", x"60", x"7C", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"60", x"60", x"7C", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"60", x"6E", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"66", x"66", x"66", x"7E", x"66", x"66", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"06", x"06", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"6C", x"78", x"70", x"78", x"6C", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"42", x"66", x"7E", x"66", x"66", x"66", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"46", x"66", x"76", x"7E", x"6E", x"66", x"62", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"66", x"66", x"7C", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"66", x"66", x"6E", x"6E", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"66", x"66", x"7C", x"78", x"6C", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"60", x"3C", x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"66", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"66", x"66", x"3C", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"7E", x"7E", x"66", x"42", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"66", x"66", x"3C", x"18", x"3C", x"66", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"06", x"0C", x"18", x"30", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"64", x"5C", x"5C", x"64", x"38", x"00", x"00", x"38", x"64", x"5C", x"5C", x"64", x"38", x"00", x"00", x"00", x"65", x"96", x"94", x"94", x"64", x"00", x"00", x"00", x"65", x"96", x"94", x"94", x"64", x"00", x"00", x"10", x"30", x"7F", x"FF", x"00", x"00", x"00", x"00", x"10", x"30", x"7F", x"FF", x"00", x"00", x"00", x"00", x"08", x"0C", x"FE", x"FF", x"00", x"00", x"00", x"00", x"08", x"0C", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"88", x"88", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"88", x"88", x"FF", x"00", x"00", x"00", x"00", x"00", 
															x"42", x"42", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"42", x"42", x"FF", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"10", x"10", x"FF", x"00", x"00", x"00", x"00", x"00", x"84", x"84", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"84", x"84", x"FF", x"00", x"00", x"00", x"00", x"00", x"21", x"21", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"21", x"21", x"FF", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"08", x"08", x"FF", x"00", x"00", x"00", x"00", x"00", x"5F", x"5F", x"DF", x"00", x"F7", x"F7", x"F7", x"00", x"40", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"88", x"88", x"FF", x"00", x"00", x"00", x"00", x"00", x"88", x"88", x"FF", x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"FF", x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"FF", x"00", x"00", x"00", x"00", x"00", 
															x"10", x"10", x"FF", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"FF", x"00", x"00", x"00", x"00", x"00", x"84", x"84", x"FF", x"00", x"00", x"00", x"00", x"00", x"84", x"84", x"FF", x"00", x"00", x"00", x"00", x"00", x"21", x"21", x"FF", x"00", x"00", x"00", x"00", x"00", x"21", x"21", x"FF", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"FF", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"FF", x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"43", x"06", x"08", x"10", x"20", x"40", x"80", x"00", x"00", x"06", x"0E", x"1C", x"38", x"70", x"E0", x"C0", x"80", x"04", x"08", x"04", x"10", x"20", x"40", x"00", x"00", x"B7", x"16", x"18", x"2E", x"52", x"A1", x"C2", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"34", x"37", x"33", x"3E", x"36", x"33", x"3F", x"20", x"2F", x"2F", x"2C", x"2F", x"2B", x"2F", x"00", x"00", x"50", x"10", x"10", x"00", x"10", x"10", x"FC", x"04", x"A4", x"E4", x"04", x"74", x"44", x"C4", x"33", x"3E", x"3C", x"17", x"13", x"0C", x"0F", x"07", x"2C", x"2D", x"37", x"1B", x"1E", x"0B", x"0C", x"07", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"24", x"64", x"44", x"A8", x"68", x"D0", x"10", x"E0", x"00", x"40", x"E0", x"90", x"80", x"82", x"82", x"81", x"07", x"5F", x"E0", x"9F", x"88", x"8A", x"8A", x"88", x"00", x"02", x"07", x"09", x"01", x"01", x"01", x"81", x"E0", x"FA", x"07", x"F9", x"11", x"11", x"11", x"11", x"86", x"87", x"83", x"40", x"30", x"08", x"18", x"00", x"94", x"94", x"90", x"49", x"37", x"08", x"1F", x"03", 
															x"81", x"C1", x"81", x"02", x"0C", x"10", x"18", x"00", x"09", x"09", x"09", x"92", x"EC", x"10", x"F8", x"C0", x"00", x"03", x"03", x"03", x"3F", x"3F", x"01", x"03", x"00", x"03", x"02", x"02", x"3E", x"20", x"3E", x"02", x"00", x"C0", x"80", x"80", x"BC", x"F8", x"80", x"80", x"00", x"C0", x"40", x"40", x"7C", x"04", x"7C", x"40", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"03", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"C0", x"00", x"03", x"63", x"30", x"3F", x"10", x"30", x"20", x"03", x"07", x"67", x"37", x"3F", x"13", x"33", x"20", x"00", x"C0", x"40", x"40", x"E0", x"80", x"80", x"00", x"C0", x"20", x"A6", x"AC", x"FC", x"48", x"4C", x"04", x"2F", x"2F", x"2F", x"4F", x"48", x"40", x"40", x"35", x"2F", x"2F", x"2F", x"5F", x"5F", x"5F", x"40", x"3F", 
															x"E0", x"E0", x"A0", x"F0", x"F0", x"00", x"00", x"00", x"F4", x"D4", x"D4", x"CA", x"0A", x"FA", x"02", x"FC", x"00", x"00", x"03", x"03", x"01", x"41", x"23", x"27", x"00", x"00", x"00", x"03", x"01", x"41", x"23", x"27", x"00", x"00", x"C0", x"C0", x"00", x"06", x"C0", x"00", x"00", x"00", x"00", x"E0", x"C0", x"C6", x"F5", x"F9", x"26", x"26", x"26", x"1F", x"07", x"01", x"02", x"00", x"27", x"3F", x"3F", x"1F", x"07", x"01", x"03", x"0F", x"00", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"F9", x"F9", x"F9", x"F6", x"E0", x"80", x"C0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"1A", x"20", x"28", x"30", x"38", x"40", x"80", x"00", x"1A", x"25", x"3E", x"25", x"35", x"6E", x"C0", x"80", x"02", x"04", x"08", x"10", x"20", x"40", x"80", x"00", x"03", x"06", x"0C", x"1E", x"34", x"60", x"F0", x"20", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"2F", x"77", x"FB", x"FD", x"FE", x"80", x"0F", x"1F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"E0", x"10", x"08", x"14", x"22", x"40", x"80", x"FF", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"FF", x"FF", x"00", x"7E", x"3D", x"1B", x"07", x"07", x"00", x"00", x"FF", x"FF", x"FF", x"7F", x"3F", x"1F", x"0F", x"00", x"FF", x"80", x"40", x"20", x"10", x"08", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"00", x"07", x"1C", x"3F", x"3F", x"3F", x"2F", x"19", x"07", x"00", x"03", x"08", x"00", x"20", x"30", x"1E", x"07", x"E0", x"F8", x"FC", x"FC", x"F8", x"E8", x"60", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"78", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"10", x"20", x"20", x"20", x"10", x"18", x"07", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"08", x"04", x"04", x"04", x"08", x"18", x"E0", x"03", x"04", x"0A", x"16", x"2E", x"3C", x"38", x"38", x"03", x"07", x"0F", x"1F", x"3F", x"3F", x"3F", x"3F", x"80", x"00", x"40", x"20", x"10", x"08", x"08", x"08", x"C0", x"E0", x"F0", x"F8", x"FC", x"FC", x"FC", x"FC", x"38", x"38", x"38", x"3C", x"16", x"0B", x"04", x"03", x"3F", x"3F", x"3F", x"3F", x"1F", x"0F", x"07", x"03", x"08", x"00", x"00", x"10", x"20", x"40", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"F8", x"F0", x"E0", x"C0", x"7F", x"7F", x"7F", x"00", x"F7", x"FF", x"80", x"BD", x"00", x"00", x"00", x"00", x"00", x"FF", x"80", x"BD", x"7F", x"7F", x"7F", x"00", x"F7", x"FF", x"00", x"EC", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"EC", x"7F", x"7F", x"7F", x"00", x"F7", x"FF", x"00", x"37", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"37", 
															x"7F", x"7F", x"7F", x"40", x"DF", x"DF", x"07", x"C7", x"00", x"00", x"7F", x"40", x"5F", x"DF", x"07", x"C7", x"7F", x"7F", x"F7", x"11", x"D1", x"D0", x"00", x"7B", x"0C", x"0E", x"F7", x"12", x"D6", x"DD", x"1B", x"7F", x"7F", x"5F", x"FF", x"C0", x"F7", x"77", x"30", x"E3", x"30", x"50", x"E0", x"40", x"60", x"F7", x"30", x"E3", x"7F", x"7F", x"7F", x"00", x"F7", x"F7", x"0F", x"F4", x"00", x"00", x"00", x"00", x"00", x"F0", x"08", x"F4", x"BD", x"98", x"58", x"5F", x"5F", x"58", x"98", x"BD", x"BD", x"98", x"58", x"5F", x"5F", x"58", x"98", x"BD", x"EC", x"C6", x"C7", x"C3", x"C1", x"C1", x"C1", x"E3", x"EC", x"C6", x"C7", x"C3", x"C1", x"C1", x"C1", x"E3", x"37", x"63", x"E3", x"C3", x"83", x"83", x"83", x"C7", x"37", x"63", x"E3", x"C3", x"83", x"83", x"83", x"C7", x"E7", x"77", x"36", x"36", x"36", x"36", x"76", x"E7", x"E7", x"77", x"37", x"37", x"36", x"3F", x"7F", x"F7",
															x"7B", x"31", x"31", x"31", x"31", x"31", x"31", x"7B", x"7F", x"F9", x"B1", x"71", x"F1", x"B1", x"31", x"7B", x"F3", x"B9", x"99", x"99", x"99", x"99", x"B9", x"F3", x"F3", x"B9", x"99", x"99", x"99", x"99", x"B9", x"F3", x"FB", x"99", x"A3", x"E4", x"E7", x"A3", x"99", x"FA", x"FA", x"99", x"A2", x"E4", x"E4", x"A2", x"99", x"FA", x"BD", x"80", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"BD", x"80", x"FF", x"00", x"00", x"00", x"00", x"00", x"E3", x"00", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"E3", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"C7", x"00", x"FE", x"00", x"F0", x"F0", x"F0", x"01", x"C7", x"00", x"FF", x"03", x"06", x"0D", x"0B", x"0F", x"C7", x"07", x"07", x"0F", x"1F", x"3F", x"00", x"FF", x"EF", x"DF", x"B7", x"6F", x"DF", x"BF", x"00", x"FF", x"7B", x"00", x"03", x"07", x"FE", x"FC", x"01", x"FF", x"7B", x"00", x"03", x"07", x"FE", x"FC", x"01", x"FF", 
															x"E3", x"00", x"3F", x"40", x"F7", x"F7", x"F7", x"00", x"E3", x"00", x"3F", x"40", x"80", x"80", x"00", x"00", x"02", x"04", x"01", x"07", x"0F", x"0F", x"1E", x"30", x"00", x"01", x"06", x"0E", x"1C", x"10", x"20", x"00", x"00", x"0F", x"81", x"01", x"C0", x"F8", x"FC", x"9F", x"60", x"8C", x"02", x"02", x"01", x"01", x"01", x"20", x"00", x"00", x"C0", x"30", x"C8", x"F4", x"F4", x"FA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"1C", x"6B", x"49", x"20", x"00", x"00", x"18", x"2C", x"2B", x"48", x"48", x"20", x"00", x"00", x"3F", x"7F", x"E7", x"C6", x"0F", x"0F", x"07", x"03", x"40", x"80", x"00", x"00", x"00", x"10", x"08", x"04", x"FA", x"FD", x"7D", x"7D", x"3D", x"3D", x"1D", x"1D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"08", x"04", x"08", x"91", x"D1", x"11", x"21", x"21", x"10", x"08", x"10", x"E1", x"91", 
															x"1D", x"D9", x"D1", x"D1", x"22", x"42", x"E4", x"20", x"00", x"00", x"00", x"00", x"80", x"80", x"20", x"20", x"00", x"00", x"07", x"19", x"E4", x"48", x"80", x"00", x"00", x"07", x"08", x"20", x"84", x"48", x"80", x"00", x"BB", x"9F", x"DF", x"BE", x"F9", x"71", x"D5", x"B4", x"FF", x"F8", x"F0", x"F0", x"E1", x"E1", x"E5", x"F4", x"5B", x"F5", x"FF", x"07", x"63", x"48", x"4A", x"02", x"0F", x"00", x"00", x"00", x"60", x"48", x"4A", x"02", x"BB", x"9D", x"94", x"E4", x"F5", x"FB", x"FC", x"7D", x"FF", x"FF", x"3F", x"0F", x"07", x"07", x"01", x"01", x"B0", x"92", x"D2", x"BA", x"EC", x"6F", x"DF", x"BD", x"F0", x"F2", x"E2", x"E2", x"F0", x"F8", x"FC", x"FE", x"40", x"48", x"48", x"6D", x"FD", x"8F", x"FF", x"FF", x"40", x"48", x"48", x"6D", x"05", x"00", x"00", x"00", x"7D", x"73", x"62", x"63", x"66", x"BD", x"DE", x"FE", x"01", x"08", x"10", x"00", x"00", x"00", x"00", x"00", 
															x"FE", x"7F", x"9E", x"1F", x"FE", x"7F", x"CE", x"4F", x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"20", x"3F", x"9F", x"57", x"BF", x"76", x"FD", x"AB", x"50", x"40", x"60", x"28", x"40", x"09", x"82", x"D0", x"F8", x"FC", x"7D", x"F2", x"7D", x"F0", x"58", x"D0", x"05", x"00", x"02", x"08", x"00", x"05", x"20", x"55", x"A7", x"B3", x"89", x"84", x"84", x"C2", x"61", x"F8", x"8C", x"BF", x"8F", x"87", x"87", x"C3", x"F1", x"F8", x"FC", x"5B", x"A5", x"14", x"1A", x"91", x"13", x"12", x"09", x"7F", x"BF", x"1F", x"1F", x"9F", x"9F", x"1F", x"0F", x"00", x"80", x"C0", x"B4", x"C9", x"6B", x"DE", x"BD", x"44", x"80", x"E0", x"FE", x"FF", x"FF", x"FF", x"FF", x"09", x"0D", x"05", x"02", x"E0", x"61", x"90", x"BA", x"0F", x"0F", x"07", x"03", x"E1", x"E1", x"F1", x"FE", x"C5", x"82", x"C1", x"A1", x"C1", x"20", x"88", x"84", x"C7", x"E3", x"E1", x"E1", x"F1", x"B8", x"8C", x"84", 
															x"93", x"89", x"C4", x"84", x"C9", x"8B", x"16", x"15", x"DF", x"EF", x"C7", x"C7", x"CF", x"8F", x"1F", x"1F", x"C0", x"B0", x"CC", x"B5", x"E9", x"6B", x"DC", x"BD", x"C0", x"F0", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"1B", x"15", x"08", x"04", x"85", x"05", x"C0", x"B2", x"1F", x"1F", x"0F", x"07", x"87", x"87", x"C7", x"FB", x"00", x"41", x"80", x"40", x"84", x"40", x"08", x"40", x"00", x"40", x"23", x"9E", x"7A", x"04", x"08", x"40", x"38", x"C4", x"3B", x"44", x"01", x"10", x"40", x"00", x"00", x"38", x"C4", x"03", x"06", x"18", x"40", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"00", x"00", x"00", x"00", x"F0", x"F0", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"10", x"F0", x"F0", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"FF", x"FF", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"7F", x"FF", x"30", x"30", x"30", x"30", x"30", x"30", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"30", x"30", x"30", x"30", x"70", x"E0", x"C0", x"80", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"80", x"30", x"30", x"30", x"30", x"3F", x"3F", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"FF", x"FF", 
															x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BF", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"F7", x"0F", x"FF", x"00", x"F7", x"F7", x"F7", x"00", x"F4", x"08", x"F0", x"00", x"00", x"00", x"00", x"00", x"EA", x"4E", x"4A", x"4A", x"4A", x"00", x"00", x"00", x"EA", x"4E", x"4A", x"4A", x"4A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00");
	
	constant ICE_CLIMBER_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"13", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"11", x"0D", x"0B", x"1B", x"1F", x"3D", x"1C", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1B", x"17", x"37", x"3F", x"7F", x"0F", x"0E", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"70", x"F8", x"F8", x"FC", x"E4", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"0F", x"1E", x"1C", x"3F", x"3F", x"38", x"00", x"00", x"00", x"01", x"03", x"00", x"00", x"07", x"78", x"7C", x"FF", x"FF", x"37", x"03", x"00", x"00", x"07", x"03", x"C0", x"F0", x"30", x"00", x"00", x"00", 
															x"C0", x"F8", x"F0", x"FC", x"FE", x"9C", x"BE", x"FE", x"00", x"00", x"00", x"00", x"00", x"60", x"40", x"00", x"7C", x"74", x"FC", x"D8", x"78", x"F0", x"F8", x"7C", x"80", x"88", x"00", x"20", x"80", x"00", x"78", x"7C", x"1C", x"3A", x"71", x"E1", x"C3", x"C6", x"6C", x"38", x"00", x"06", x"0F", x"1F", x"3F", x"3E", x"1C", x"18", x"06", x"09", x"13", x"26", x"4C", x"98", x"B0", x"60", x"00", x"07", x"0F", x"1E", x"3C", x"78", x"70", x"60", x"4E", x"2C", x"18", x"00", x"00", x"00", x"00", x"00", x"34", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"0C", x"0C", x"0C", x"06", x"06", x"46", x"3C", x"78", x"30", x"10", x"30", x"78", x"7C", x"78", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"43", x"43", x"67", x"26", x"2A", x"22", x"16", x"14", x"FC", x"FC", x"F8", x"78", x"74", x"7C", x"38", x"38", x"3C", x"1C", x"18", x"08", x"00", x"00", x"00", x"00", x"38", x"18", x"10", x"00", x"00", x"00", x"00", x"00", x"26", x"12", x"01", x"41", x"08", x"01", x"04", x"00", x"11", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"30", x"00", x"04", x"20", x"10", x"00", x"00", x"10", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"44", x"00", x"00", x"20", x"04", x"00", x"00", x"02", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"01", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"3A", x"5C", x"BE", x"5F", x"3E", x"1C", x"00", x"01", x"3A", x"5C", x"BE", x"5F", x"3E", x"1C", x"00", x"18", x"3C", x"7E", x"5F", x"2D", x"32", x"4C", x"80", x"18", x"3C", x"7E", x"5F", x"2D", x"32", x"4C", x"80", 
															x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"1A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"03", x"07", x"0E", x"07", x"01", x"03", x"07", x"0F", x"1C", x"08", x"00", x"00", x"01", x"03", x"00", x"00", x"0F", x"1F", x"1E", x"1D", x"3B", x"3B", x"03", x"81", x"00", x"00", x"00", x"00", x"00", x"04", x"3D", x"3F", x"C0", x"E0", x"F0", x"7C", x"7E", x"38", x"10", x"00", x"1F", x"9F", x"8F", x"47", x"6E", x"38", x"10", x"00", x"00", x"00", x"4C", x"FC", x"FC", x"78", x"08", x"7C", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"7C", x"DC", x"FC", x"F8", x"F8", x"FC", x"FC", x"BC", x"00", x"04", x"04", x"08", x"C0", x"00", x"00", x"04", x"7C", x"7C", x"F8", x"F8", x"F8", x"F0", x"82", x"3A", x"0C", x"0C", x"18", x"38", x"70", x"EC", x"FC", x"CC", x"7C", x"7C", x"FE", x"FE", x"7E", x"1E", x"3C", x"78", x"8C", x"8C", x"06", x"06", x"02", x"02", x"04", x"00", 
															x"00", x"00", x"00", x"01", x"02", x"02", x"1A", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"1C", x"07", x"0E", x"07", x"01", x"03", x"07", x"0F", x"0F", x"08", x"00", x"00", x"01", x"03", x"00", x"00", x"00", x"1F", x"1F", x"1F", x"3F", x"3C", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"03", x"3F", x"3F", x"1E", x"01", x"03", x"03", x"0F", x"1F", x"00", x"01", x"03", x"1E", x"0C", x"04", x"02", x"01", x"00", x"00", x"00", x"00", x"4C", x"FC", x"FC", x"78", x"08", x"7C", x"7C", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"DC", x"FC", x"F8", x"FC", x"FC", x"FE", x"FE", x"DE", x"04", x"04", x"08", x"C0", x"00", x"00", x"02", x"02", x"DE", x"DE", x"DC", x"BC", x"38", x"7A", x"72", x"B8", x"02", x"06", x"04", x"0C", x"8C", x"1C", x"1C", x"3C", x"FC", x"FC", x"F8", x"F8", x"F0", x"F8", x"F8", x"E0", x"0C", x"1C", x"18", x"38", x"30", x"18", x"18", x"20", 
															x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"1A", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"03", x"07", x"0E", x"07", x"01", x"03", x"07", x"0F", x"1C", x"08", x"00", x"00", x"01", x"03", x"00", x"00", x"0F", x"1F", x"1F", x"1F", x"3F", x"3E", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"01", x"3F", x"3C", x"07", x"0F", x"0F", x"0F", x"3F", x"7F", x"1F", x"07", x"18", x"10", x"00", x"00", x"01", x"01", x"1B", x"07", x"00", x"00", x"4C", x"FC", x"FC", x"78", x"08", x"7C", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"7C", x"DC", x"FC", x"F8", x"FC", x"FE", x"FE", x"FE", x"00", x"04", x"04", x"08", x"C0", x"00", x"02", x"02", x"EF", x"EF", x"F7", x"F7", x"F7", x"07", x"0F", x"8B", x"03", x"03", x"13", x"31", x"31", x"F1", x"E1", x"61", x"C6", x"E0", x"E7", x"EF", x"BF", x"9F", x"06", x"06", x"3A", x"7C", x"FF", x"F3", x"81", x"81", x"02", x"02", 
															x"7E", x"FE", x"C0", x"CE", x"C6", x"FE", x"7E", x"00", x"01", x"01", x"3F", x"21", x"29", x"01", x"81", x"7F", x"7C", x"FE", x"C6", x"C6", x"C6", x"FE", x"7C", x"00", x"02", x"01", x"39", x"21", x"21", x"01", x"83", x"7E", x"38", x"7C", x"EE", x"C6", x"FE", x"FE", x"C6", x"00", x"04", x"02", x"11", x"29", x"01", x"01", x"39", x"C7", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"21", x"21", x"21", x"11", x"83", x"46", x"2C", x"18", x"6C", x"FE", x"FE", x"D6", x"D6", x"D6", x"C6", x"00", x"12", x"01", x"01", x"29", x"29", x"29", x"39", x"E7", x"7E", x"FE", x"C0", x"FC", x"C0", x"FE", x"7E", x"00", x"01", x"01", x"3F", x"02", x"3E", x"01", x"81", x"7F", x"70", x"98", x"68", x"78", x"D8", x"78", x"F8", x"70", x"0C", x"06", x"67", x"77", x"D7", x"77", x"06", x"0C", x"7C", x"FE", x"C6", x"DE", x"DC", x"CE", x"C6", x"00", x"02", x"01", x"39", x"21", x"22", x"31", x"29", x"E7", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"1F", x"0F", x"1F", x"3F", x"3D", x"00", x"01", x"01", x"01", x"10", x"20", x"07", x"0D", x"3F", x"7F", x"7F", x"31", x"00", x"04", x"04", x"08", x"00", x"00", x"1E", x"3E", x"0F", x"0B", x"1B", x"17", x"3F", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"F0", x"E0", x"F0", x"F8", x"78", x"F0", x"E0", x"E0", x"C0", x"10", x"08", x"C0", x"60", x"C0", x"F0", x"F8", x"F8", x"80", x"40", x"4C", x"28", x"00", x"00", x"F0", x"F8", x"EC", x"AC", x"BC", x"D8", x"F8", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"01", x"07", x"0E", x"1F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"70", x"F0", x"F0", x"E0", x"00", x"00", x"38", x"FE", x"9E", x"1C", x"3C", x"FE", x"FF", x"00", x"00", x"02", x"01", x"00", x"00", x"00", x"00", x"1F", x"3F", x"31", x"60", x"C0", x"80", x"00", x"00", x"00", x"00", x"03", x"1F", x"1F", x"0F", x"0F", x"0F", x"1F", x"3F", x"3C", x"60", x"60", x"30", x"30", x"70", x"1F", x"3F", x"FF", x"FF", x"FF", x"7F", x"3F", x"34", x"E0", x"C0", x"00", x"00", x"01", x"1D", x"3F", x"34", x"00", x"00", x"C0", x"FE", x"F0", x"C0", x"80", x"80", x"C0", x"F8", x"3E", x"01", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"E0", x"80", x"00", x"00", x"47", x"2E", x"1C", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"01", x"07", x"0E", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"78", x"C0", x"03", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"70", x"F0", x"F0", x"E0", x"00", x"00", x"38", x"FE", x"9E", x"1C", x"3C", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"1F", x"FF", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"3F", x"20", x"1E", x"1F", x"BF", x"7F", x"3F", x"3C", x"34", x"DF", x"E1", x"E0", x"40", x"01", x"1F", x"3C", x"34", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"F0", x"FC", x"00", x"00", x"E0", x"F0", x"C0", x"00", x"00", x"00", x"FF", x"FC", x"10", x"0E", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"34", x"FF", x"FF", x"FF", x"7F", x"3F", x"1F", x"3F", x"35", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"81", x"00", x"40", x"20", x"10", x"00", x"00", x"00", x"00", x"E7", x"BE", x"DC", x"EF", x"F0", x"FF", x"FE", x"F8", x"01", x"03", x"03", x"07", x"01", x"00", x"00", x"06", x"01", x"03", x"03", x"07", x"03", x"07", x"07", x"09", x"04", x"00", x"10", x"30", x"20", x"00", x"00", x"00", x"19", x"3F", x"6F", x"4F", x"5F", x"7F", x"3F", x"1F", x"E0", x"F0", x"F0", x"F0", x"B8", x"80", x"00", x"C0", x"E0", x"F0", x"F0", x"F0", x"F8", x"F0", x"F0", x"30", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"F0", x"F0", x"F0", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"0E", x"1F", x"13", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"11", x"0D", x"0B", x"1B", x"1D", x"3D", x"1C", x"0F", x"00", x"0C", x"0A", x"1A", x"1E", x"00", x"0C", x"1F", 
															x"1B", x"17", x"37", x"3E", x"0E", x"00", x"0E", x"1E", x"1B", x"17", x"37", x"3F", x"7F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"60", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"70", x"70", x"70", x"70", x"70", x"60", x"C0", x"60", x"80", x"00", x"80", x"E8", x"7C", x"04", x"00", x"00", x"E0", x"70", x"F8", x"F0", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"09", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"05", x"0D", x"0E", x"1E", x"0E", x"00", x"0B", x"06", x"05", x"0D", x"0F", x"00", x"00", x"0F", x"07", x"14", x"15", x"05", x"07", x"07", x"0F", x"00", x"01", x"0C", x"0D", x"3D", x"3F", x"1F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"C0", x"60", x"30", x"38", 
															x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"80", x"38", x"38", x"38", x"38", x"30", x"60", x"30", x"B8", x"C0", x"D8", x"FC", x"C0", x"C0", x"80", x"E0", x"E0", x"D8", x"D8", x"FC", x"F8", x"FC", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"09", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"05", x"0D", x"0E", x"1E", x"6E", x"60", x"08", x"06", x"05", x"0D", x"0F", x"00", x"60", x"7F", x"3F", x"00", x"11", x"02", x"71", x"38", x"18", x"00", x"00", x"3F", x"0F", x"3E", x"0F", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"C0", x"60", x"30", x"38", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"02", x"4C", x"38", x"38", x"38", x"38", x"30", x"60", x"3A", x"7C", x"EC", x"70", x"F8", x"78", x"B6", x"6E", x"06", x"0E", x"FC", x"78", x"FE", x"7C", x"B8", x"F0", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"30", x"79", x"3F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"0F", x"2F", x"BB", x"E7", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0E", x"07", x"07", x"03", x"03", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"FE", x"DE", x"E7", x"D7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"9B", x"E7", x"AF", x"FF", x"FE", x"FC", x"7E", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6F", x"47", x"E7", x"F2", x"C0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"71", x"7D", x"7F", x"00", x"00", x"00", x"00", x"3E", x"71", x"7D", x"7F", x"08", x"14", x"2A", x"5E", x"7E", x"7C", x"3A", x"11", x"08", x"14", x"2A", x"5E", x"7E", x"7C", x"3A", x"11", 
															x"01", x"00", x"00", x"00", x"00", x"00", x"03", x"02", x"01", x"00", x"00", x"00", x"03", x"07", x"04", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"17", x"3E", x"3B", x"6E", x"FC", x"F0", x"A4", x"EE", x"6E", x"7C", x"7C", x"38", x"00", x"00", x"A4", x"EE", x"6E", x"7C", x"FC", x"F8", x"E0", x"F0", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"03", x"02", x"06", x"07", x"0F", x"07", x"00", x"00", x"03", x"02", x"06", x"07", x"00", x"01", x"0C", x"06", x"1A", x"0B", x"03", x"01", x"6E", x"37", x"1B", x"1A", x"1E", x"07", x"1F", x"3F", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"00", x"00", x"00", x"00", x"00", x"60", x"30", x"18", 
															x"60", x"60", x"E0", x"E0", x"60", x"60", x"00", x"00", x"1C", x"1C", x"9C", x"9C", x"9C", x"18", x"30", x"00", x"E0", x"FE", x"EC", x"E0", x"C0", x"01", x"04", x"C0", x"FC", x"FE", x"FC", x"F8", x"F8", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"07", x"0F", x"00", x"10", x"00", x"00", x"01", x"01", x"00", x"00", x"1F", x"0F", x"00", x"20", x"00", x"00", x"00", x"01", x"03", x"07", x"3E", x"1E", x"7F", x"7F", x"FF", x"06", x"00", x"00", x"7F", x"3E", x"08", x"08", x"E8", x"F8", x"3C", x"1C", x"7F", x"3E", x"08", x"08", x"08", x"0C", x"0A", x"1B", x"DC", x"A4", x"A4", x"C4", x"84", x"88", x"00", x"00", x"DB", x"BB", x"BB", x"FB", x"3A", x"34", x"30", x"20", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"80", x"60", x"40", x"C0", x"E0", x"80", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"0E", x"1F", x"13", x"11", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"ED", x"EB", x"43", x"01", x"00", x"00", x"00", x"00", x"EC", x"FA", x"7A", x"3E", x"1F", x"0F", x"0F", x"07", x"0A", x"01", x"09", x"00", x"01", x"05", x"07", x"03", x"05", x"0E", x"06", x"0F", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"80", x"C0", x"60", x"70", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"70", x"70", x"70", x"70", x"60", x"C0", x"E0", x"F0", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"80", x"F0", x"F8", x"78", x"FC", x"F8", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"03", x"9C", x"8C", x"6C", x"5C", x"DC", x"EC", x"68", x"20", x"03", x"03", x"63", x"53", x"D3", x"F3", x"67", x"00", 
															x"00", x"00", x"00", x"64", x"76", x"5F", x"8F", x"86", x"1F", x"3D", x"38", x"72", x"61", x"40", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"60", x"70", x"F8", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"03", x"04", x"00", x"08", x"00", x"00", x"00", x"00", x"04", x"03", x"07", x"06", x"0E", x"1F", x"0F", x"00", x"00", x"01", x"00", x"01", x"00", x"00", x"00", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"78", x"5C", x"8C", x"EC", x"DC", x"93", x"E3", x"00", x"04", x"02", x"02", x"E3", x"D3", x"9F", x"FF", 
															x"C2", x"04", x"00", x"00", x"00", x"00", x"00", x"06", x"3E", x"FA", x"B8", x"70", x"70", x"78", x"FC", x"F8", x"0E", x"8E", x"C2", x"C0", x"80", x"00", x"00", x"00", x"E0", x"70", x"20", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"02", x"00", x"00", x"08", x"11", x"01", x"01", x"03", x"03", x"01", x"01", x"01", x"01", x"3B", x"12", x"40", x"70", x"60", x"60", x"00", x"00", x"04", x"0D", x"0E", x"0E", x"1E", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B0", x"F8", x"5C", x"0C", x"2C", x"1C", x"1C", x"08", x"80", x"84", x"82", x"82", x"E3", x"D3", x"F3", x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F6", x"FE", x"F8", x"F0", x"70", x"70", x"F0", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"04", x"3C", x"FE", x"F1", x"43", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"43", x"E3", x"FF", x"F3", x"E3", x"67", x"3F", x"7F", x"0C", x"1C", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"F7", x"F7", x"F7", x"FB", x"7E", x"F8", x"A8", x"10", x"30", x"30", x"10", x"18", x"0D", x"0B", x"0F", x"20", x"00", x"30", x"3F", x"1F", x"1F", x"03", x"07", x"47", x"3F", x"0F", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"DC", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C4", x"FF", x"FE", x"FF", x"FE", x"F2", x"F0", x"E0", x"F0", x"43", x"40", x"40", x"58", x"90", x"F0", x"E0", x"70", x"F0", x"F8", x"F0", x"EC", x"9D", x"3F", x"3F", x"3F", x"30", x"38", x"18", x"1C", x"64", x"C4", x"C1", x"C1", x"3F", x"1F", x"0E", x"06", x"C0", x"C0", x"80", x"00", x"C3", x"E3", x"82", x"02", x"C0", x"40", x"00", x"00", 
															x"00", x"1D", x"0F", x"3F", x"10", x"34", x"31", x"1F", x"00", x"00", x"00", x"00", x"0F", x"0B", x"CE", x"E0", x"1F", x"3F", x"3F", x"3F", x"1F", x"1F", x"2B", x"7E", x"60", x"00", x"03", x"07", x"06", x"00", x"34", x"7E", x"00", x"C0", x"F0", x"F8", x"DC", x"E8", x"FC", x"FA", x"00", x"00", x"00", x"00", x"20", x"10", x"00", x"04", x"FE", x"F4", x"FA", x"FF", x"ED", x"FB", x"5E", x"0C", x"60", x"E8", x"E4", x"C1", x"13", x"07", x"0E", x"0C", x"0E", x"07", x"1F", x"08", x"1A", x"18", x"0F", x"0F", x"00", x"00", x"00", x"07", x"05", x"67", x"70", x"30", x"1F", x"1F", x"1F", x"0F", x"0F", x"05", x"0E", x"01", x"00", x"00", x"00", x"00", x"00", x"02", x"0E", x"01", x"E0", x"F8", x"FC", x"6E", x"74", x"FE", x"FD", x"FF", x"00", x"00", x"00", x"90", x"88", x"00", x"02", x"30", x"FA", x"FD", x"FF", x"F6", x"FC", x"B8", x"C0", x"F0", x"3C", x"1A", x"38", x"38", x"00", x"40", x"F0", x"F0", 
															x"0E", x"07", x"1F", x"08", x"1A", x"18", x"0F", x"0F", x"00", x"00", x"00", x"07", x"05", x"67", x"70", x"30", x"1F", x"1F", x"1F", x"6F", x"2F", x"35", x"18", x"00", x"00", x"00", x"00", x"70", x"30", x"38", x"18", x"00", x"E0", x"F8", x"FC", x"6E", x"74", x"FE", x"FD", x"FF", x"00", x"00", x"00", x"90", x"88", x"00", x"02", x"30", x"FE", x"FF", x"FF", x"F6", x"FC", x"B2", x"1E", x"3C", x"3C", x"1E", x"06", x"0E", x"00", x"0E", x"1E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"30", x"38", x"58", x"58", x"DC", x"DC", x"9C", x"BE", x"08", x"04", x"26", x"26", x"32", x"32", x"6B", x"41", x"00", x"00", x"3D", x"7C", x"78", x"F3", x"E2", x"60", x"00", x"00", x"3D", x"7F", x"7F", x"FC", x"FC", x"7F", x"27", x"2F", x"16", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"3F", x"1F", x"1F", x"0F", x"03", 
															x"00", x"70", x"F8", x"1C", x"04", x"61", x"23", x"06", x"00", x"70", x"F8", x"FC", x"FC", x"9D", x"9F", x"FF", x"CC", x"E8", x"70", x"10", x"08", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"E0", x"00", x"00", x"01", x"33", x"73", x"0A", x"02", x"47", x"00", x"38", x"7D", x"4F", x"0F", x"06", x"0E", x"59", x"6F", x"6F", x"2F", x"1F", x"0F", x"07", x"03", x"03", x"71", x"70", x"30", x"00", x"10", x"08", x"35", x"13", x"00", x"70", x"D0", x"F0", x"EC", x"FC", x"34", x"3C", x"00", x"00", x"00", x"08", x"90", x"E0", x"20", x"20", x"30", x"98", x"F0", x"80", x"B8", x"08", x"08", x"C8", x"38", x"98", x"7C", x"7E", x"46", x"C6", x"86", x"C4", x"01", x"03", x"07", x"07", x"07", x"07", x"05", x"07", x"01", x"03", x"07", x"07", x"05", x"05", x"05", x"07", x"06", x"0F", x"1B", x"3F", x"55", x"7F", x"6E", x"3C", x"07", x"0F", x"1F", x"3F", x"7F", x"7F", x"7E", x"3C", 
															x"80", x"C0", x"E0", x"E0", x"E0", x"E0", x"60", x"E0", x"80", x"C0", x"E0", x"E0", x"60", x"60", x"60", x"E0", x"C0", x"C0", x"40", x"80", x"80", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"03", x"07", x"07", x"0F", x"0F", x"0F", x"0F", x"01", x"11", x"3B", x"5F", x"0F", x"0F", x"07", x"01", x"0F", x"0E", x"0E", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"00", x"40", x"00", x"60", x"00", x"80", x"C0", x"E0", x"E0", x"F0", x"F0", x"F0", x"F0", x"60", x"88", x"DC", x"FA", x"F0", x"F0", x"E0", x"80", x"F0", x"70", x"30", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"06", x"16", x"06", x"00", x"03", x"07", x"1F", x"3D", x"39", x"7B", x"7B", x"7F", x"00", x"10", x"01", x"00", x"08", x"00", x"00", x"00", x"7F", x"7F", x"3F", x"3F", x"3F", x"3F", x"1F", x"07", 
															x"00", x"00", x"00", x"80", x"C0", x"C0", x"D0", x"00", x"C0", x"E0", x"F0", x"78", x"38", x"BC", x"BC", x"FC", x"00", x"08", x"00", x"20", x"00", x"80", x"00", x"00", x"FC", x"FC", x"FC", x"F8", x"F8", x"F0", x"E0", x"C0", x"06", x"07", x"03", x"01", x"01", x"01", x"03", x"03", x"06", x"07", x"03", x"01", x"01", x"01", x"03", x"03", x"0F", x"1F", x"1D", x"1D", x"1F", x"0E", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"60", x"60", x"40", x"D8", x"B8", x"E0", x"80", x"20", x"60", x"60", x"40", x"D8", x"B8", x"E0", x"80", x"E0", x"F0", x"70", x"70", x"F0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"13", x"26", x"6C", x"4C", x"48", x"48", x"00", x"01", x"1B", x"3F", x"7F", x"7D", x"79", x"79", x"4C", x"4C", x"44", x"44", x"20", x"24", x"16", x"1A", x"7F", x"7F", x"7F", x"7C", x"30", x"3F", x"1F", x"1B", 
															x"00", x"00", x"98", x"10", x"08", x"08", x"08", x"08", x"80", x"80", x"DC", x"FE", x"FE", x"BE", x"9E", x"9E", x"08", x"08", x"10", x"10", x"00", x"10", x"10", x"00", x"FE", x"FC", x"FC", x"3C", x"0C", x"F8", x"F8", x"D0", x"05", x"0F", x"17", x"3F", x"1F", x"1F", x"1F", x"0F", x"05", x"0F", x"17", x"3E", x"1E", x"1A", x"1C", x"0E", x"0F", x"0F", x"1F", x"1D", x"19", x"1F", x"1E", x"0F", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"B0", x"F8", x"F8", x"F0", x"E8", x"F0", x"E0", x"20", x"B0", x"F8", x"F8", x"B0", x"68", x"F0", x"60", x"E0", x"E0", x"F0", x"70", x"30", x"F0", x"F0", x"E0", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"11", x"0D", x"0B", x"1B", x"1D", x"3F", x"1F", x"00", x"00", x"0C", x"0A", x"1A", x"1E", x"00", x"00", x"1F", x"10", x"00", x"2C", x"0C", x"00", x"00", x"0E", x"1E", x"0F", x"1D", x"1F", x"3F", x"7C", x"0F", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"70", x"70", x"70", x"70", x"70", x"60", x"C0", x"E0", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"E0", x"F0", x"B8", x"70", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"05", x"0D", x"0E", x"1F", x"0F", x"00", x"08", x"06", x"05", x"0D", x"0F", x"00", x"00", x"0F", x"07", x"10", x"10", x"00", x"00", x"00", x"0E", x"00", x"01", x"1F", x"0B", x"39", x"3D", x"1F", x"01", x"00", x"00", x"88", x"5C", x"3E", x"7E", x"7A", x"54", x"28", x"10", x"88", x"5C", x"3E", x"7E", x"7A", x"54", x"28", x"10", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"00", x"00", x"38", x"38", x"38", x"38", x"30", x"60", x"F0", x"B0", 
															x"00", x"00", x"C0", x"C0", x"00", x"00", x"E0", x"E0", x"B8", x"78", x"E8", x"D8", x"FC", x"F0", x"00", x"00", x"14", x"15", x"05", x"07", x"07", x"03", x"0C", x"1D", x"0C", x"0D", x"3D", x"3F", x"1F", x"0F", x"00", x"00", x"06", x"05", x"0D", x"0E", x"1F", x"6F", x"60", x"08", x"06", x"05", x"0D", x"0F", x"00", x"60", x"7F", x"37", x"00", x"10", x"00", x"70", x"38", x"18", x"00", x"00", x"3F", x"0E", x"3E", x"0F", x"07", x"01", x"00", x"00", x"0C", x"1E", x"3F", x"3E", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"23", x"1F", x"0E", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"00", x"00", x"38", x"38", x"38", x"38", x"30", x"60", x"F8", x"FC", x"0C", x"0C", x"00", x"00", x"06", x"0E", x"06", x"0C", x"DC", x"EC", x"7E", x"3C", x"F8", x"F0", x"00", x"00", x"00", x"20", x"30", x"00", x"00", x"00", x"0C", x"1D", x"1D", x"3D", x"2C", x"1E", x"3E", x"0F", x"00", x"00", 
															x"00", x"00", x"F0", x"F8", x"78", x"18", x"1C", x"0C", x"38", x"7C", x"0E", x"06", x"06", x"06", x"03", x"83", x"0C", x"0C", x"2E", x"3E", x"3F", x"7F", x"3F", x"18", x"B3", x"73", x"D1", x"01", x"00", x"60", x"30", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"38", x"00", x"00", x"00", x"00", x"00", x"E0", x"E0", x"C0", x"28", x"2C", x"1E", x"7E", x"3F", x"80", x"80", x"00", x"C0", x"C4", x"EE", x"FE", x"FF", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"83", x"BF", x"00", x"20", x"31", x"21", x"61", x"01", x"00", x"00", x"7F", x"DF", x"0E", x"1E", x"7E", x"3E", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"10", x"38", x"28", x"00", x"00", x"00", x"00", x"E0", x"E0", x"C0", x"C0", x"2C", x"1E", x"7E", x"3F", x"80", x"80", x"80", x"00", x"C4", x"EE", x"FE", x"FF", x"60", x"00", x"00", x"00", 
															x"00", x"80", x"00", x"04", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"00", x"00", x"0F", x"3F", x"3F", x"00", x"01", x"01", x"1F", x"1F", x"10", x"00", x"0F", x"3F", x"7F", x"7F", x"01", x"04", x"04", x"08", x"00", x"00", x"1E", x"3E", x"31", x"0B", x"1B", x"17", x"3F", x"0E", x"00", x"00", x"00", x"10", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"00", x"00", x"E0", x"F8", x"F8", x"F0", x"E0", x"E0", x"F0", x"F0", x"10", x"00", x"C0", x"C0", x"F8", x"F8", x"C0", x"40", x"4C", x"28", x"00", x"00", x"F0", x"F8", x"EC", x"AC", x"BC", x"D8", x"F8", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"00", x"00", x"00", x"00", x"00", x"0F", x"10", x"20", x"1D", x"3D", x"3F", x"3B", x"3C", x"3F", x"1F", x"0F", x"25", x"0D", x"1F", x"1B", x"1C", x"0F", x"07", x"30", 
															x"01", x"04", x"04", x"68", x"20", x"00", x"1E", x"3E", x"7E", x"7B", x"6B", x"77", x"3F", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"00", x"00", x"00", x"00", x"00", x"E0", x"10", x"08", x"70", x"78", x"F8", x"B8", x"78", x"F8", x"F0", x"E0", x"48", x"60", x"F0", x"B0", x"70", x"E0", x"C0", x"18", x"00", x"40", x"40", x"2C", x"09", x"03", x"F3", x"FA", x"FC", x"BC", x"AC", x"DC", x"FC", x"E4", x"04", x"04", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"0F", x"1F", x"DD", x"FD", x"FF", x"33", x"30", x"0F", x"10", x"20", x"E5", x"CD", x"DF", x"D0", x"D0", x"38", x"1F", x"6F", x"E1", x"E4", x"E8", x"E0", x"40", x"48", x"27", x"10", x"1E", x"1B", x"17", x"1F", x"37", x"00", x"C0", x"F8", x"F8", x"F8", x"F8", x"F8", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"E0", x"F0", x"73", x"7B", x"FB", x"98", x"18", x"E2", x"12", x"0A", x"4B", x"63", x"F3", x"17", x"16", x"38", x"F0", x"EC", x"0E", x"4E", x"2E", x"0E", x"04", x"24", x"C8", x"10", x"F0", x"B0", x"D0", x"F0", x"D8", x"07", x"0F", x"1F", x"1F", x"3D", x"3F", x"3F", x"1F", x"07", x"0F", x"1D", x"1D", x"3D", x"3F", x"3F", x"1F", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"00", x"03", x"07", x"07", x"0F", x"1F", x"1E", x"1D", x"0F", x"E0", x"F0", x"F8", x"F8", x"7C", x"FC", x"FC", x"F8", x"E0", x"F0", x"78", x"78", x"7C", x"FC", x"FC", x"F8", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"40", x"40", x"80", x"80", x"00", x"60", x"F0", x"F8", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"18", x"F0", x"E0", x"00", x"7C", x"FE", x"FF", x"FD", x"FC", x"78", x"00", x"00", x"00", x"00", x"00", x"02", x"03", x"87", x"FE", x"7C", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"23", x"E0", x"60", x"AA", x"23", x"E8", x"48", x"50", x"23", x"F0", x"48", x"AF", x"20", x"62", x"01", x"77", x"20", x"63", x"5A", x"7A", x"20", x"7D", x"01", x"7C", x"20", x"82", x"C9", x"78", x"21", x"A2", x"01", x"79", x"21", x"A3", x"5A", x"7B", x"20", x"9D", x"C9", x"7D", x"21", x"BD", x"01", x"7E", x"20", x"83", x"5A", x"FD", x"20", x"A3", x"5A", x"FD", x"20", x"C3", x"5A", x"FD", x"20", x"E3", x"5A", x"FD", x"21", x"03", x"5A", x"FD", x"20", x"8B", x"0A", x"5E", x"FD", x"FD", x"60", x"61", x"61", x"FD", x"60", x"61", x"61", x"20", x"AB", x"0A", x"5F", x"FD", x"FD", x"5F", x"62", x"FD", x"FD", x"5F", x"66", x"68", x"20", x"CB", x"0A", x"5F", x"FD", x"FD", 
															x"5F", x"63", x"FD", x"FD", x"5F", x"67", x"69", x"20", x"EB", x"0A", x"5F", x"FD", x"FD", x"64", x"65", x"61", x"FD", x"64", x"65", x"61", x"21", x"23", x"1A", x"60", x"61", x"61", x"FD", x"5E", x"FD", x"FD", x"FD", x"5E", x"FD", x"60", x"6A", x"60", x"6A", x"FD", x"60", x"61", x"6A", x"FD", x"60", x"61", x"61", x"FD", x"60", x"61", x"6A", x"21", x"43", x"1A", x"5F", x"62", x"FD", x"FD", x"5F", x"FD", x"FD", x"FD", x"5F", x"FD", x"5F", x"6B", x"6C", x"6D", x"FD", x"5F", x"6E", x"71", x"FD", x"5F", x"66", x"68", x"FD", x"5F", x"6E", x"71", x"21", x"63", x"1A", x"5F", x"63", x"FD", x"FD", x"5F", x"63", x"FD", x"FD", x"5F", x"FD", x"5F", x"74", x"75", x"5F", x"FD", x"5F", x"6F", x"72", x"FD", x"5F", x"67", x"69", x"FD", x"5F", x"76", x"72", x"21", x"83", x"1A", x"64", x"65", x"61", x"FD", x"64", x"65", x"61", x"FD", x"5F", x"FD", x"5F", x"FD", x"FD", x"5F", x"FD", x"5F", x"70", x"73", 
															x"FD", x"64", x"65", x"61", x"FD", x"5F", x"FD", x"5F", x"22", x"0A", x"0D", x"01", x"38", x"8D", x"37", x"33", x"A3", x"3D", x"8E", x"38", x"36", x"33", x"3C", x"3D", x"22", x"4A", x"0D", x"02", x"38", x"8D", x"37", x"33", x"A3", x"3D", x"8E", x"38", x"36", x"33", x"3C", x"3D", x"22", x"8A", x"08", x"3C", x"5B", x"93", x"5A", x"3A", x"33", x"3B", x"5A", x"22", x"CA", x"03", x"7F", x"80", x"81", x"22", x"D2", x"05", x"00", x"3E", x"3F", x"40", x"41", x"23", x"05", x"01", x"83", x"23", x"0B", x"05", x"00", x"3E", x"3F", x"40", x"41", x"23", x"12", x"02", x"82", x"83", x"23", x"19", x"05", x"00", x"3E", x"3F", x"40", x"41", x"23", x"69", x"0E", x"FC", x"01", x"09", x"08", x"04", x"38", x"5A", x"3B", x"5A", x"3A", x"3D", x"5A", x"35", x"5B", x"00", x"3F", x"00", x"14", x"0F", x"31", x"12", x"30", x"0F", x"25", x"29", x"0A", x"0F", x"30", x"21", x"01", x"0F", x"27", x"17", x"07", x"0F", 
															x"30", x"12", x"26", x"00", x"23", x"CC", x"44", x"55", x"23", x"D4", x"44", x"55", x"23", x"DC", x"44", x"55", x"23", x"E4", x"44", x"55", x"23", x"EC", x"44", x"55", x"23", x"F4", x"44", x"55", x"21", x"08", x"06", x"5A", x"5B", x"38", x"38", x"38", x"38", x"21", x"28", x"06", x"34", x"5B", x"5A", x"93", x"91", x"39", x"20", x"6A", x"08", x"3C", x"5B", x"93", x"5A", x"3A", x"33", x"3B", x"5A", x"20", x"82", x"01", x"95", x"20", x"A2", x"D6", x"96", x"23", x"62", x"01", x"97", x"20", x"83", x"4C", x"98", x"23", x"63", x"4C", x"99", x"20", x"8F", x"01", x"9A", x"20", x"AF", x"D6", x"9B", x"23", x"6F", x"01", x"9C", x"20", x"C5", x"08", x"01", x"38", x"8D", x"37", x"33", x"A3", x"3D", x"8E", x"22", x"C6", x"05", x"3A", x"5B", x"3A", x"33", x"37", x"22", x"E4", x"83", x"84", x"85", x"86", x"22", x"E5", x"48", x"87", x"23", x"25", x"48", x"88", x"22", x"ED", x"83", x"89", x"8A", x"8B", 
															x"23", x"0B", x"01", x"00", x"00", x"21", x"16", x"06", x"5A", x"5B", x"38", x"38", x"38", x"38", x"21", x"36", x"06", x"34", x"5B", x"5A", x"93", x"91", x"39", x"20", x"90", x"01", x"95", x"20", x"B0", x"D6", x"96", x"23", x"70", x"01", x"97", x"20", x"91", x"4C", x"98", x"23", x"71", x"4C", x"99", x"20", x"9D", x"01", x"9A", x"20", x"BD", x"D6", x"9B", x"23", x"7D", x"01", x"9C", x"20", x"D3", x"08", x"02", x"38", x"8D", x"37", x"33", x"A3", x"3D", x"8E", x"22", x"D4", x"05", x"3A", x"5B", x"3A", x"33", x"37", x"22", x"F2", x"83", x"84", x"85", x"86", x"22", x"F3", x"48", x"87", x"23", x"33", x"48", x"88", x"22", x"FB", x"83", x"89", x"8A", x"8B", x"23", x"19", x"01", x"00", x"00", x"3F", x"00", x"08", x"0F", x"30", x"21", x"11", x"0F", x"30", x"25", x"15", x"3F", x"10", x"0C", x"0F", x"30", x"11", x"26", x"0F", x"30", x"15", x"26", x"0F", x"30", x"21", x"12", x"00", x"FF", x"FF", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"55", x"AA", x"55", x"22", x"88", x"00", x"22", x"00", x"AA", x"55", x"AA", x"DD", x"77", x"FF", x"DD", x"00", x"00", x"08", x"00", x"00", x"00", x"80", x"00", x"FF", x"FF", x"F7", x"FF", x"FF", x"FF", x"7F", x"FF", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"60", x"C0", x"DE", x"C6", x"66", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"38", x"38", x"10", x"10", x"10", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"19", x"1F", x"1F", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"BF", x"8C", x"8C", x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"3C", x"7C", x"70", x"3C", x"0E", x"7E", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E7", x"FF", x"7E", x"3C", x"3C", x"3C", x"3C", x"3C", x"00", x"0C", x"8F", x"CF", x"CF", x"CF", x"CF", x"CF", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"7E", x"FF", x"E7", x"C3", x"C3", x"C3", x"C3", x"C3", x"00", x"C0", x"F8", x"FC", x"FC", x"FC", x"FC", x"FC", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"7E", x"7E", x"66", x"66", x"7A", x"7C", x"00", x"FF", x"C1", x"A3", x"9F", x"9F", x"BB", x"FD", x"FF", 
															x"E0", x"F0", x"70", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"30", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"7E", x"FF", x"E7", x"C3", x"C3", x"C3", x"C3", x"C3", x"00", x"C0", x"F8", x"FC", x"FC", x"FC", x"FC", x"FC", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"00", x"00", x"07", x"0C", x"08", x"08", x"00", x"00", x"00", x"0F", x"18", x"10", x"10", x"10", x"07", x"0F", x"0E", x"0C", x"0C", x"0C", x"0C", x"0C", x"00", x"00", x"01", x"03", x"03", x"03", x"03", x"03", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", 
															x"7E", x"FF", x"E7", x"C3", x"C3", x"C3", x"C3", x"C3", x"00", x"03", x"1F", x"3F", x"3F", x"3F", x"3F", x"3F", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"0F", x"1F", x"19", x"11", x"11", x"13", x"1F", x"0F", x"00", x"00", x"07", x"0F", x"0F", x"0F", x"1F", x"0F", x"7F", x"FF", x"C3", x"81", x"81", x"C3", x"FF", x"7F", x"00", x"00", x"3D", x"7F", x"7F", x"7F", x"FF", x"7F", x"60", x"F0", x"D0", x"90", x"90", x"B0", x"F0", x"60", x"00", x"00", x"30", x"70", x"70", x"70", x"F0", x"60", x"0F", x"1F", x"18", x"10", x"10", x"18", x"1F", x"0F", x"00", x"00", x"07", x"0F", x"0F", x"0F", x"1F", x"0F", 
															x"EF", x"FF", x"78", x"30", x"30", x"78", x"FF", x"EF", x"00", x"00", x"A7", x"EF", x"EF", x"EF", x"FF", x"EF", x"E0", x"F0", x"30", x"10", x"10", x"30", x"F0", x"E0", x"00", x"00", x"D0", x"F0", x"F0", x"F0", x"F0", x"E0", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"42", x"24", x"18", x"18", x"24", x"42", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", 
															x"FC", x"F0", x"E0", x"C0", x"C0", x"80", x"80", x"80", x"00", x"00", x"01", x"07", x"0F", x"0F", x"1F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"C0", x"C0", x"E0", x"F0", x"FC", x"3F", x"3F", x"3F", x"1F", x"1F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"7F", x"FF", x"FF", x"E0", x"E0", x"E0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"07", x"07", x"E0", x"E0", x"E0", x"E0", x"FF", x"FF", x"7F", x"3F", x"07", x"07", x"07", x"07", x"00", x"00", x"00", x"80", 
															x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"1F", x"07", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"F0", x"FC", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"60", x"F0", x"F0", x"F0", x"F0", x"F0", x"FF", x"FF", x"9F", x"0F", x"07", x"07", x"03", x"03", x"00", x"00", x"06", x"0F", x"0F", x"0F", x"0F", x"0F", x"3F", x"BF", x"F9", x"F0", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"3F", x"3F", x"3E", x"7F", x"FF", x"FE", x"E0", x"E0", x"E0", x"E0", x"C1", x"80", x"00", x"00", x"00", x"00", x"07", x"07", x"E0", x"E0", x"E0", x"E0", x"FE", x"FF", x"FF", x"FE", x"07", x"07", x"07", x"07", x"01", x"00", x"00", x"00", 
															x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"07", x"FF", x"FF", x"7F", x"7F", x"7E", x"FE", x"FC", x"F8", x"1F", x"07", x"03", x"01", x"01", x"00", x"00", x"00", x"E0", x"E0", x"E0", x"F8", x"FC", x"FE", x"7F", x"7F", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"07", x"7F", x"FF", x"FF", x"FF", x"FE", x"FE", x"FC", x"F8", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"E0", x"E0", x"FE", x"FF", x"FF", x"FF", x"07", x"07", x"07", x"07", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"40", x"20", x"10", x"0F", x"08", x"08", x"08", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"FF", x"FF", x"FF", x"F8", x"F0", x"E0", x"C0", x"80", x"08", x"08", x"08", x"08", x"0F", x"1F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"E0", x"E0", x"00", x"01", x"03", x"07", x"FF", x"0F", x"0F", x"0F", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"F7", x"FB", x"FD", x"FE", x"FC", x"FD", x"31", x"31", x"31", x"31", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"F3", x"FB", x"9B", x"9B", x"9B", x"FB", x"F3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"30", x"F6", x"E6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"06", x"06", x"06", x"06", x"06", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"60", x"60", x"66", x"66", x"60", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0C", x"08", x"08", x"00", x"00", x"1F", x"30", x"20", x"20", x"20", x"20", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"08", x"0C", x"07", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"30", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"60", x"20", x"20", x"00", x"00", x"F0", x"18", x"08", x"08", x"08", x"08", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"20", x"60", x"C0", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"18", x"F0", x"00", x"00", x"00", x"00", x"3A", x"5C", x"66", x"66", x"3A", x"5C", x"00", x"77", x"81", x"81", x"9A", x"1F", x"9B", x"9D", x"EE", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5C", x"3A", x"66", x"66", x"5C", x"3A", x"00", x"EE", x"81", x"83", x"1F", x"9E", x"9D", x"BB", x"77", 
															x"7F", x"FF", x"C3", x"81", x"81", x"C3", x"FF", x"7F", x"00", x"00", x"3D", x"7F", x"7F", x"7F", x"FF", x"7F", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"C1", x"C1", x"7F", x"00", x"00", x"00", x"00", x"00", x"3F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"D6", x"FE", x"FE", x"EE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"38", x"70", x"60", x"60", x"60", x"00", x"0F", x"1F", x"38", x"73", x"67", x"6E", x"6C", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"61", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"60", x"60", x"60", x"70", x"38", x"1F", x"0F", x"00", x"6C", x"6E", x"67", x"73", x"38", x"1F", x"0F", x"00", 
															x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"F0", x"F8", x"1C", x"0E", x"06", x"06", x"06", x"00", x"F0", x"F8", x"1C", x"CE", x"E6", x"76", x"36", x"86", x"86", x"86", x"86", x"86", x"86", x"86", x"86", x"36", x"36", x"36", x"36", x"36", x"36", x"36", x"36", x"06", x"06", x"06", x"0E", x"1C", x"F8", x"F0", x"00", x"36", x"76", x"E6", x"CE", x"1C", x"F8", x"F0", x"00", x"E7", x"FF", x"7E", x"3C", x"3C", x"3C", x"3C", x"3C", x"00", x"30", x"F1", x"F3", x"F3", x"F3", x"F3", x"F3", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"3C", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"7E", x"FF", x"E7", x"C3", x"C3", x"C3", x"C3", x"C3", x"00", x"03", x"1F", x"3F", x"3F", x"3F", x"3F", x"3F", 
															x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"C3", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"00", x"7E", x"7E", x"66", x"66", x"7A", x"7C", x"00", x"FF", x"C1", x"A3", x"9F", x"9F", x"BB", x"FD", x"FF", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"40", x"20", x"08", x"50", x"20", x"30", x"04", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"42", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0A", x"01", x"20", x"14", x"81", x"04", x"28", x"54", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"AA", x"55", x"AA", x"55", x"AA", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"C0", x"60", x"20", x"20", x"00", x"00", x"00", x"E0", x"30", x"10", x"10", x"10", x"00", x"38", x"0C", x"4C", x"86", x"06", x"4B", x"01", x"FF", x"C7", x"F3", x"F3", x"F9", x"F9", x"F4", x"FE", x"00", x"00", x"00", x"08", x"20", x"00", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"38", x"5C", x"5C", x"8E", x"4A", x"86", x"26", x"FF", x"C7", x"E3", x"E3", x"F1", x"F5", x"F9", x"F9", x"82", x"12", x"42", x"01", x"10", x"81", x"0A", x"45", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"8A", x"55", x"AA", x"55", x"AA", x"D5", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", 
															x"00", x"00", x"00", x"40", x"60", x"24", x"1A", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"0B", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"02", x"15", x"0E", x"05", x"02", x"14", x"01", x"2A", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"04", x"80", x"48", x"80", x"40", x"A8", x"54", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AA", x"55", x"AA", x"57", x"BF", x"5F", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1C", x"7E", x"DE", x"0F", x"9F", x"07", x"A3", x"00", x"E3", x"81", x"21", x"F0", x"E0", x"F8", x"FC", x"FF", 
															x"80", x"20", x"80", x"00", x"40", x"80", x"00", x"20", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"04", x"00", x"00", x"40", x"00", x"80", x"21", x"50", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A1", x"52", x"A9", x"53", x"BD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"08", x"0C", x"07", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"18", x"0F", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"60", x"60", x"70", x"38", x"3C", x"00", x"00", x"00", x"80", x"80", x"80", x"C0", x"C0", x"7C", x"FC", x"CC", x"86", x"06", x"82", x"83", x"C3", x"80", x"00", x"30", x"78", x"F8", x"7C", x"7C", x"3C", x"C3", x"47", x"47", x"47", x"43", x"42", x"04", x"00", x"3C", x"B8", x"B8", x"B8", x"BC", x"BD", x"FB", x"FF", x"00", x"00", x"20", x"1A", x"04", x"80", x"40", x"A0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"50", x"EA", x"75", x"AA", x"F5", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"60", x"30", x"38", x"18", x"0C", x"1C", x"7C", x"9C", x"80", x"C0", x"C0", x"E0", x"F0", x"E0", x"80", x"60", x"0E", x"0E", x"06", x"26", x"D2", x"EA", x"F7", x"FF", x"F0", x"F0", x"F8", x"F8", x"FC", x"FC", x"FE", x"FE", x"20", x"60", x"C0", x"00", x"00", x"00", x"00", x"00", x"10", x"10", x"30", x"E0", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"03", x"02", x"06", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"07", x"07", x"07", x"07", x"07", x"0E", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"03", x"1D", x"1C", x"18", x"1D", x"3A", x"35", x"7F", x"FF", x"03", x"03", x"07", x"07", x"0F", x"1F", x"3F", x"7F", x"EE", x"DD", x"00", x"00", x"00", x"DD", x"BB", x"00", x"00", x"00", x"BB", x"77", x"EE", x"DD", x"BB", x"77", x"01", x"01", x"03", x"07", x"06", x"0E", x"0C", x"08", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"07", x"18", x"38", x"30", x"32", x"74", x"7C", x"7C", x"7C", x"07", x"07", x"0F", x"0D", x"0B", x"03", x"03", x"03", 
															x"DC", x"D8", x"88", x"08", x"08", x"01", x"21", x"41", x"23", x"27", x"77", x"F7", x"F7", x"FE", x"FE", x"FE", x"01", x"03", x"02", x"82", x"C2", x"20", x"01", x"02", x"FE", x"FC", x"FD", x"7D", x"3D", x"DF", x"FF", x"FF", x"05", x"12", x"A9", x"57", x"BF", x"77", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"77", x"BB", x"00", x"00", x"00", x"BB", x"DD", x"00", x"00", x"00", x"DD", x"EE", x"77", x"BB", x"DD", x"EE", x"00", x"04", x"00", x"00", x"20", x"00", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"04", x"08", x"08", x"10", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"38", x"70", x"E2", x"E6", x"C2", x"81", x"81", x"FF", x"C7", x"8F", x"1F", x"1F", x"3F", x"7F", x"7F", x"02", x"01", x"04", x"01", x"0A", x"81", x"4A", x"A4", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"57", x"AE", x"D7", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"04", x"00", x"40", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"04", x"00", x"00", x"20", x"00", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"02", x"24", x"18", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"84", x"00", x"80", x"01", x"A0", x"02", x"45", x"8A", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"55", x"AA", x"D4", x"A9", x"D2", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"20", x"02", x"00", x"00", x"08", x"00", x"40", x"00", x"00", x"02", x"00", x"00", x"00", x"02", x"00", x"00", 
															x"00", x"06", x"1F", x"1D", x"3C", x"38", x"39", x"30", x"FF", x"F9", x"E0", x"E2", x"C3", x"C7", x"C7", x"CF", x"31", x"30", x"78", x"78", x"68", x"C0", x"81", x"80", x"CF", x"CF", x"87", x"87", x"97", x"3F", x"7F", x"7F", x"00", x"04", x"00", x"00", x"20", x"00", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"02", x"84", x"00", x"21", x"00", x"48", x"22", x"45", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"2A", x"55", x"AA", x"75", x"BB", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"02", x"40", x"01", x"00", x"00", x"00", x"80", x"08", x"00", x"40", x"01", x"10", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"80", x"44", x"80", x"40", x"C0", x"FF", x"FF", x"FF", x"7F", x"FF", x"FF", x"FF", x"FF", x"20", x"50", x"24", x"90", x"00", x"24", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"10", x"02", x"20", x"04", x"51", x"22", x"54", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AA", x"55", x"AA", x"75", x"BA", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7E", x"7E", x"66", x"66", x"7A", x"7C", x"00", x"FF", x"C1", x"A3", x"9F", x"9F", x"BB", x"FD", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"38", x"38", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"3C", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"66", x"06", x"1E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"70", x"60", x"7E", x"7E", x"7E", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"66", x"06", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"06", x"66", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"1C", x"3C", x"3C", x"6C", x"6C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6C", x"7E", x"7E", x"7E", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"60", x"7C", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"66", x"7E", x"7E", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"66", x"60", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"66", x"66", x"7E", x"7E", x"3C", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"66", x"0E", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"66", x"66", x"7E", x"7E", x"3C", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF");
	
	constant ROAD_FIGHTER_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F9", x"F9", x"F9", x"F9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F3", x"F3", x"F3", x"F3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"E7", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CF", x"CF", x"CF", x"CF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"9F", x"9F", x"9F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"CF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"0F", x"6F", x"6F", x"6F", x"6F", x"6F", x"6F", x"0F", x"8F", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"8F", x"FC", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"1F", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"1F", x"1F", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"1F", x"F8", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"F8", x"06", x"03", x"03", x"03", x"03", x"03", x"03", x"06", 
															x"3F", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"3F", x"3F", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"3F", x"F0", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"F0", x"0C", x"07", x"07", x"07", x"07", x"07", x"07", x"0C", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"E0", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"E0", x"18", x"0E", x"0E", x"0E", x"0E", x"0E", x"0E", x"18", x"C1", x"ED", x"ED", x"ED", x"ED", x"ED", x"ED", x"C1", x"31", x"1D", x"1D", x"1D", x"1D", x"1D", x"1D", x"31", x"83", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"83", x"63", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"63", x"07", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"07", x"C7", x"77", x"77", x"77", x"77", x"77", x"77", x"C7", x"1F", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"1F", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"80", 
															x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"3F", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"F8", x"FE", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FE", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F0", x"FC", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"FC", x"E1", x"ED", x"ED", x"ED", x"ED", x"ED", x"ED", x"E1", x"F8", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F8", x"C3", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"C3", x"F0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"F0", x"87", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"87", x"E0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"E0", 
															x"0F", x"6F", x"6F", x"6F", x"6F", x"6F", x"6F", x"0F", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"C0", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"05", x"0B", x"17", x"5F", x"3F", x"3F", x"FF", x"FD", x"FF", x"F4", x"F8", x"F0", x"E0", x"C0", x"80", x"08", x"41", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"7F", x"3F", x"1F", x"0F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"1F", x"1F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"1F", x"1F", x"41", x"10", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"13", x"43", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"7F", x"FF", x"7F", x"7F", x"7F", x"FF", x"7F", x"7F", x"80", x"80", x"80", x"80", x"80", x"A0", x"B8", x"BC", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0F", x"07", x"07", x"03", x"00", x"07", x"0F", x"1F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"FC", x"FC", x"00", x"FC", x"FC", x"FC", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7F", x"7F", x"7E", x"7E", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"BF", x"BF", x"3F", x"FC", x"FC", x"00", x"FC", x"FC", x"3C", x"BC", x"3C", x"FC", x"FC", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"7F", x"7E", x"7E", x"7F", x"7F", x"7F", x"7F", x"00", x"FF", x"BF", x"BF", x"3F", x"FF", x"FF", x"FF", x"03", x"FC", x"3C", x"BC", x"3C", x"FC", x"FC", x"FC", x"00", x"7E", x"7D", x"7A", x"75", x"6A", x"55", x"2A", x"55", x"BE", x"BD", x"BA", x"B5", x"AA", x"95", x"AA", x"95", x"BF", x"5F", x"AF", x"57", x"AA", x"54", x"AA", x"54", x"BF", x"5F", x"AF", x"57", x"AA", x"54", x"AA", x"54", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"00", x"00", x"00", x"00", x"6A", x"35", x"1A", x"25", x"0A", x"11", x"06", x"01", x"AA", x"D5", x"EA", x"FD", x"F6", x"EF", x"FB", x"FF", x"A8", x"50", x"A8", x"50", x"A0", x"50", x"A0", x"72", x"A8", x"50", x"A8", x"50", x"A0", x"50", x"50", x"DF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"0B", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"7F", x"7F", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"0F", x"1F", x"FF", x"FF", x"00", x"00", x"01", x"07", x"0F", x"1F", x"00", x"00", x"0F", x"7E", x"FD", x"FE", x"FD", x"FA", x"FF", x"FF", x"0F", x"7E", x"FD", x"FE", x"FD", x"FA", x"C2", x"A8", x"70", x"B2", x"58", x"AD", x"52", x"AA", x"3D", x"57", x"0F", x"8D", x"47", x"A2", x"55", x"A9", x"E0", x"E0", x"E1", x"E3", x"E3", x"E3", x"E3", x"E3", x"60", x"60", x"61", x"63", x"60", x"63", x"63", x"63", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"7F", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", 
															x"FD", x"FA", x"F5", x"FA", x"F5", x"FA", x"FD", x"FE", x"FD", x"FA", x"F5", x"FA", x"05", x"F2", x"F9", x"FE", x"56", x"AB", x"54", x"A9", x"50", x"A1", x"40", x"80", x"55", x"AA", x"55", x"A8", x"51", x"A0", x"41", x"81", x"E3", x"E3", x"E3", x"E3", x"E3", x"E3", x"03", x"03", x"63", x"63", x"63", x"63", x"63", x"63", x"03", x"03", x"FF", x"FF", x"FF", x"DF", x"DF", x"1F", x"FF", x"FF", x"00", x"FF", x"FF", x"1F", x"5F", x"1F", x"FF", x"FF", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"1F", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"E3", x"E3", x"E3", x"E3", x"E3", x"E3", x"E3", x"E0", x"63", x"63", x"63", x"63", x"63", x"63", x"63", x"60", x"FF", x"DF", x"DF", x"1F", x"FF", x"FF", x"FF", x"00", x"FF", x"1F", x"5F", x"1F", x"FF", x"FF", x"FF", x"00", 
															x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DE", x"1C", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DE", x"1C", x"E3", x"E3", x"E3", x"E3", x"E3", x"E1", x"00", x"00", x"63", x"63", x"63", x"63", x"63", x"61", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"DB", x"6D", x"36", x"FF", x"FF", x"FF", x"FF", x"00", x"DB", x"6D", x"36", x"FC", x"F8", x"F0", x"E0", x"00", x"60", x"B0", x"D8", x"FC", x"F8", x"F0", x"E0", x"00", x"60", x"B0", x"D8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"7F", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"FC", x"F8", x"FF", x"FF", x"FF", x"FF", x"F1", x"FF", x"FF", x"F9", x"FF", x"FF", x"7F", x"97", x"17", x"8B", x"07", x"17", x"FF", x"7F", x"EF", x"5F", x"DF", x"57", x"FF", x"AB", 
															x"E0", x"C3", x"C4", x"88", x"82", x"C3", x"8F", x"FF", x"E0", x"C2", x"C3", x"8D", x"83", x"C3", x"8F", x"FF", x"04", x"21", x"03", x"29", x"47", x"57", x"7F", x"FF", x"D4", x"D1", x"7B", x"95", x"1B", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9D", x"8C", x"CD", x"C0", x"00", x"FF", x"FF", x"FF", x"9D", x"8C", x"CD", x"C0", x"00", x"01", x"C0", x"C8", x"CC", x"DC", x"9D", x"BF", x"FF", x"01", x"C0", x"C8", x"CC", x"DC", x"9D", x"BF", x"FF", x"E9", x"DA", x"F1", x"E9", x"F5", x"F2", x"E4", x"F2", x"FE", x"F5", x"DE", x"F6", x"FA", x"FD", x"FB", x"ED", x"E7", x"EA", x"C1", x"D7", x"C6", x"BB", x"5D", x"2F", x"F8", x"F5", x"FE", x"E8", x"F9", x"C4", x"A2", x"D0", x"FF", x"EF", x"FF", x"BF", x"FB", x"FF", x"EF", x"FE", x"00", x"10", x"00", x"40", x"04", x"00", x"10", x"01", x"00", x"48", x"00", x"01", x"08", x"00", x"20", x"00", x"FF", x"B7", x"FF", x"FE", x"F7", x"FF", x"DF", x"FF", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F1", x"FB", x"F3", x"F7", x"C1", x"EF", x"FD", x"FF", x"FE", x"FC", x"FE", x"EC", x"FE", x"F0", x"F5", x"E9", x"F5", x"E2", x"EB", x"E9", x"DE", x"D5", x"CA", x"F6", x"FA", x"FD", x"F4", x"D6", x"F9", x"EE", x"6F", x"F7", x"AF", x"5D", x"FF", x"77", x"FF", x"7E", x"90", x"08", x"50", x"A2", x"00", x"88", x"00", x"81", x"CD", x"A7", x"D6", x"C3", x"9D", x"CB", x"CF", x"E7", x"F2", x"F8", x"F9", x"FC", x"E2", x"F4", x"F8", x"F9", x"E1", x"F3", x"F9", x"E3", x"F8", x"F9", x"FD", x"FE", x"FE", x"FC", x"F6", x"FC", x"FF", x"FE", x"FE", x"FF", x"7F", x"FB", x"7F", x"F5", x"5F", x"FF", x"9F", x"57", x"90", x"04", x"80", x"0A", x"A0", x"02", x"60", x"A8", x"37", x"8D", x"D7", x"CD", x"CF", x"E2", x"E3", x"E5", x"C8", x"F2", x"F8", x"F2", x"F8", x"FD", x"FC", x"FE", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"64", x"94", x"84", x"87", x"84", x"84", x"94", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"9E", x"90", x"90", x"9C", x"90", x"90", x"90", x"9E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"64", x"95", x"85", x"86", x"85", x"85", x"94", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"87", x"84", x"04", x"04", x"07", x"84", x"84", x"84", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"19", x"A4", x"A4", x"A4", x"24", x"24", x"24", x"19", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D2", x"9A", x"9A", x"96", x"96", x"92", x"92", x"D2", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"FF", x"4F", x"4F", x"4F", x"4F", x"4F", x"4F", x"4F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"3F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"0F", x"1F", x"FF", x"FF", x"FF", x"FF", x"1F", x"00", x"0F", x"1F", x"FF", x"FF", x"FF", x"FF", x"1F", x"CF", x"CF", x"CF", x"CF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", x"43", x"0B", x"03", x"03", x"13", x"00", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"03", x"13", x"03", x"07", x"43", x"0B", x"03", x"23", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"00", 
															x"67", x"EF", x"D7", x"CB", x"E7", x"EF", x"B7", x"F7", x"27", x"6F", x"5E", x"4D", x"27", x"6F", x"56", x"17", x"6B", x"9C", x"AF", x"97", x"EB", x"EE", x"E3", x"F3", x"6F", x"94", x"AC", x"51", x"6B", x"2E", x"12", x"1B", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"17", x"BF", x"EF", x"E5", x"C5", x"EF", x"FF", x"83", x"07", x"B5", x"ED", x"E1", x"C1", x"EC", x"FF", x"FF", x"FF", x"FB", x"E3", x"A1", x"F7", x"FF", x"FF", x"00", x"00", x"C0", x"60", x"20", x"20", x"40", x"00", x"F9", x"E8", x"ED", x"FF", x"FF", x"81", x"0C", x"ED", x"C1", x"E0", x"E5", x"CF", x"FF", x"F1", x"9C", x"FD", x"00", x"80", x"00", x"64", x"20", x"80", x"60", x"50", x"FF", x"7F", x"FF", x"BB", x"DF", x"7F", x"DF", x"AF", 
															x"3F", x"3D", x"3E", x"7D", x"BB", x"7C", x"FA", x"FF", x"F8", x"EB", x"F5", x"E3", x"F4", x"EB", x"FD", x"EA", x"F6", x"FD", x"FF", x"FF", x"FB", x"F7", x"DF", x"FF", x"0F", x"97", x"0B", x"B0", x"84", x"89", x"6B", x"C7", x"01", x"07", x"0F", x"1E", x"3F", x"3C", x"34", x"7B", x"FF", x"FF", x"FF", x"FE", x"FD", x"FC", x"F6", x"EF", x"D0", x"F0", x"60", x"C8", x"B8", x"44", x"02", x"54", x"FF", x"FF", x"67", x"CB", x"BB", x"E7", x"C3", x"F4", x"00", x"00", x"00", x"14", x"00", x"00", x"00", x"00", x"FF", x"FF", x"E7", x"D4", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"2F", x"13", x"07", x"01", x"00", x"28", x"95", x"DC", x"6E", x"EF", x"EA", x"88", x"FF", x"FF", x"BF", x"DC", x"4E", x"EB", x"BA", x"88", x"00", x"10", x"E8", x"B0", x"D4", x"6C", x"FA", x"D4", x"FF", x"FF", x"FF", x"B3", x"D4", x"CC", x"FA", x"F4", 
															x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"30", x"30", x"70", x"70", x"70", x"70", x"70", x"70", x"30", x"30", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"FC", x"FC", x"FC", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BF", x"2F", x"27", x"7F", x"EF", x"C5", x"E5", x"EF", x"A7", x"1F", x"07", x"65", x"ED", x"C3", x"E1", x"EC", x"FD", x"F1", x"D8", x"F5", x"FD", x"FF", x"FF", x"FF", x"FD", x"81", x"C8", x"E5", x"DD", x"FF", x"FF", x"FF", x"E7", x"E3", x"F2", x"F9", x"FC", x"FF", x"FE", x"FE", x"F9", x"FC", x"FD", x"FE", x"FF", x"FC", x"FF", x"FF", x"2D", x"4F", x"3E", x"5A", x"9F", x"36", x"BE", x"1E", x"FA", x"FD", x"FD", x"F5", x"F2", x"E9", x"F3", x"F5", 
															x"7E", x"7D", x"FA", x"FB", x"F7", x"FD", x"FF", x"EF", x"C1", x"E3", x"C5", x"95", x"8A", x"07", x"87", x"DB", x"FF", x"7B", x"BF", x"9F", x"FF", x"DC", x"D7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3B", x"37", x"09", x"1E", x"14", x"14", x"07", x"01", x"DE", x"EB", x"ED", x"FE", x"F2", x"FD", x"FF", x"FF", x"38", x"54", x"84", x"70", x"C0", x"20", x"D0", x"A0", x"F8", x"D7", x"A5", x"73", x"C7", x"6B", x"DF", x"FF", x"00", x"00", x"00", x"00", x"08", x"05", x"00", x"00", x"00", x"00", x"00", x"80", x"88", x"C5", x"DA", x"FF", x"00", x"00", x"08", x"20", x"00", x"00", x"00", x"00", x"00", x"01", x"0B", x"27", x"1B", x"AF", x"FF", x"FF", x"70", x"EA", x"78", x"E8", x"24", x"72", x"78", x"74", x"F4", x"6A", x"F8", x"AC", x"F4", x"F2", x"F8", x"D4", x"00", x"00", x"40", x"00", x"00", x"00", x"40", x"00", x"7F", x"3F", x"7F", x"3F", x"3F", x"3F", x"7F", x"7F", 
															x"70", x"EB", x"7C", x"E9", x"6F", x"7D", x"3E", x"07", x"D4", x"69", x"FC", x"AC", x"DF", x"BD", x"EE", x"FF", x"00", x"00", x"04", x"84", x"2C", x"2C", x"E9", x"ED", x"3F", x"5F", x"2D", x"84", x"4E", x"EB", x"BB", x"ED", x"F8", x"E7", x"CF", x"9F", x"BB", x"3D", x"7E", x"78", x"FF", x"F8", x"F0", x"E0", x"C4", x"CE", x"83", x"87", x"1F", x"E7", x"F3", x"F9", x"FD", x"8C", x"7E", x"7E", x"FF", x"1F", x"0F", x"47", x"83", x"F3", x"B1", x"89", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FB", x"EB", x"EB", x"FB", x"FF", x"FF", x"FF", x"FF", x"38", x"28", x"28", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"3F", x"3F", x"1F", x"1F", x"0F", x"0F", x"F9", x"F9", x"F9", x"F9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"07", x"07", x"0F", x"3F", x"3F", x"7F", x"7F", x"FF", x"5F", x"2F", x"5E", x"B6", x"BD", x"6B", x"57", x"CF", x"5F", x"AF", x"46", x"8F", x"FF", x"FF", x"FF", x"F9", x"FF", x"1F", x"FF", x"F8", x"F0", x"00", x"C0", x"E6", x"F8", x"E2", x"8F", x"97", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7E", x"0C", x"00", x"00", x"03", x"FF", x"FF", x"FF", x"BF", x"7F", x"FF", x"FC", x"E3", x"FF", x"FF", x"F0", x"C0", x"80", x"1F", x"3F", x"9C", x"80", x"60", x"FF", x"FD", x"FA", x"DE", x"7C", x"DC", x"B0", x"E0", x"87", x"3F", x"34", x"3A", x"84", x"34", x"48", x"30", x"00", x"00", x"02", x"04", x"04", x"08", x"08", x"10", x"03", x"03", x"03", x"03", x"07", x"07", x"0F", x"1F", x"7F", x"7F", x"FF", x"37", x"3F", x"5F", x"2F", x"1B", x"47", x"6F", x"F9", x"A7", x"BF", x"DE", x"EF", x"FB", 
															x"3C", x"68", x"3C", x"18", x"00", x"00", x"00", x"00", x"FC", x"E8", x"DC", x"E9", x"FF", x"FF", x"FF", x"FF", x"BB", x"19", x"10", x"10", x"EC", x"CE", x"8C", x"89", x"C3", x"E5", x"EE", x"EE", x"12", x"30", x"70", x"F1", x"7A", x"76", x"3E", x"BF", x"9F", x"CF", x"E7", x"F8", x"85", x"89", x"C1", x"C0", x"E0", x"F0", x"F8", x"FF", x"3E", x"DE", x"DC", x"7D", x"F9", x"F3", x"E7", x"1F", x"C1", x"21", x"23", x"83", x"07", x"0F", x"1F", x"FF", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"07", x"03", x"03", x"01", x"01", x"00", x"F3", x"F3", x"F3", x"F3", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"F8", x"E3", x"0F", x"66", x"F8", x"FF", x"F0", x"F8", x"F8", x"FC", x"FE", x"FF", x"FF", x"FF", x"00", x"80", x"C0", x"C0", x"00", x"BC", x"C3", x"62", x"10", x"08", x"00", x"04", x"04", x"01", x"02", x"02", x"0F", x"0F", x"07", x"07", x"07", x"02", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"EF", x"FB", x"ED", x"1D", x"FE", x"FF", x"05", x"0E", x"17", x"1F", x"1F", x"3F", x"6F", x"35", x"FD", x"FE", x"F6", x"D5", x"DF", x"9F", x"EF", x"85", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", 
															x"FB", x"B7", x"AF", x"9F", x"AD", x"B5", x"B9", x"FF", x"04", x"48", x"50", x"60", x"52", x"4A", x"46", x"00", x"FF", x"FF", x"FF", x"B7", x"51", x"55", x"B5", x"FF", x"00", x"00", x"00", x"48", x"AE", x"AA", x"4A", x"00", x"FF", x"FF", x"FF", x"1A", x"D8", x"1A", x"0A", x"FF", x"00", x"00", x"00", x"E5", x"27", x"E5", x"F5", x"00", x"FF", x"FF", x"EF", x"FC", x"2C", x"AC", x"AC", x"FD", x"03", x"03", x"13", x"00", x"D0", x"50", x"50", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"80", x"C0", x"40", x"20", x"00", x"00", x"00", x"80", x"00", x"00", x"80", x"80", x"80", x"80", x"FF", x"FF", x"03", x"C7", x"8F", x"87", x"FF", x"FF", x"FF", x"FF", x"03", x"C7", x"8F", x"87", x"FF", x"FF", x"FF", x"E3", x"F8", x"F8", x"F8", x"F9", x"39", x"FC", x"7F", x"FF", x"F9", x"F9", x"F9", x"F9", x"F9", x"7C", 
															x"FF", x"BF", x"4E", x"CE", x"CE", x"CE", x"8E", x"1D", x"FC", x"BE", x"CE", x"CE", x"CE", x"CE", x"8E", x"1C", x"14", x"28", x"14", x"0C", x"07", x"2F", x"56", x"B8", x"08", x"16", x"1E", x"0F", x"07", x"17", x"2E", x"78", x"00", x"7F", x"70", x"6F", x"6F", x"6F", x"6F", x"70", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"E0", x"7D", x"7D", x"FD", x"FD", x"FD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"3D", x"F8", x"FA", x"F7", x"F7", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"F8", x"FB", x"FB", x"7B", x"7B", x"BB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"1C", x"EF", x"EF", x"EF", x"EF", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"06", x"BE", x"BE", x"BE", x"BE", x"BE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"7F", x"BF", x"5F", x"AF", x"57", x"AB", x"55", x"AA", x"80", x"40", x"A0", x"50", x"A8", x"54", x"AA", x"55", x"E7", x"E7", x"E7", x"E7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FA", x"F5", x"EA", x"D5", x"AA", x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7E", x"BD", x"5A", x"A5", x"5A", x"A5", x"5A", x"00", x"80", x"40", x"A0", x"50", x"A0", x"50", x"A0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"3F", x"1F", x"1F", x"0F", x"07", x"07", x"03", x"00", x"00", x"FE", x"E0", x"E0", x"C0", x"C0", x"80", x"00", x"00", x"FE", x"E0", x"E0", x"C0", x"C0", x"80", x"FF", x"C3", x"D3", x"E9", x"E9", x"C1", x"F3", x"FF", x"00", x"30", x"30", x"18", x"18", x"38", x"30", x"00", x"3B", x"1D", x"0E", x"07", x"01", x"00", x"00", x"00", x"3B", x"1D", x"0E", x"07", x"01", x"00", x"00", x"FF", 
															x"6C", x"B6", x"DB", x"EF", x"F7", x"3B", x"0F", x"00", x"6C", x"B6", x"DB", x"EF", x"F7", x"3B", x"0F", x"FF", x"03", x"06", x"8A", x"D5", x"FE", x"C4", x"D8", x"42", x"00", x"01", x"85", x"CE", x"C3", x"BF", x"27", x"FF", x"7F", x"7F", x"7F", x"6F", x"6F", x"70", x"7F", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7D", x"7D", x"7D", x"7D", x"7D", x"FD", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EF", x"E0", x"CF", x"DF", x"DF", x"DF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B8", x"3A", x"9B", x"DB", x"DB", x"DB", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1F", x"7F", x"3F", x"9F", x"CF", x"EF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BE", x"BE", x"BE", x"BE", x"BE", x"BE", x"FE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
															x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"A5", x"5A", x"A5", x"5A", x"A5", x"5A", x"A5", x"5A", x"50", x"A0", x"50", x"A0", x"50", x"A0", x"50", x"A0", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A5", x"5A", x"A5", x"5A", x"A5", x"5A", x"BD", x"7E", x"50", x"A0", x"50", x"A0", x"50", x"A0", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"07", x"07", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"87", x"C1", x"AC", x"E6", x"F0", x"F8", x"FF", x"00", x"60", x"60", x"7C", x"3E", x"1E", x"0C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", 
															x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"6A", x"37", x"3B", x"1D", x"1A", x"0E", x"07", x"07", x"B5", x"CB", x"DE", x"E3", x"F5", x"F3", x"F9", x"FC", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"33", x"33", x"CC", x"CC", x"33", x"33", x"81", x"81", x"81", x"81", x"81", x"81", x"FF", x"FF", x"19", x"19", x"67", x"67", x"19", x"19", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"00", x"00", x"08", x"14", x"22", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"00", x"00", x"30", x"30", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CC", x"CC", x"33", x"33", x"0C", x"0C", x"33", x"33", 
															x"55", x"AA", x"55", x"AB", x"57", x"AF", x"5F", x"7F", x"AA", x"55", x"AA", x"54", x"A8", x"50", x"A0", x"80", x"55", x"AA", x"D5", x"EA", x"F5", x"FA", x"FD", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"07", x"0F", x"1F", x"1F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FD", x"DF", x"FF", x"F7", x"BF", x"FD", x"FF", x"00", x"80", x"08", x"00", x"20", x"02", x"00", x"40", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", 
															x"6C", x"F6", x"F9", x"E3", x"E7", x"9F", x"16", x"2D", x"12", x"0E", x"09", x"03", x"27", x"5C", x"96", x"25", x"80", x"40", x"00", x"00", x"00", x"00", x"40", x"80", x"7F", x"3F", x"3F", x"3F", x"3F", x"3F", x"7F", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"CD", x"CD", x"31", x"30", x"CC", x"CC", x"33", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BC", x"8C", x"8C", x"F8", x"00", x"00", x"33", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"33", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"63", x"63", x"63", x"00", x"00", x"33", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"30", x"3F", x"00", x"00", x"33", x"33", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"33", x"B3", x"0C", x"0C", x"33", x"33", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"FF", x"00", x"00", x"00", x"30", x"78", x"78", x"10", x"00", x"07", x"1F", x"BF", x"BF", x"FF", x"FF", x"FF", x"FF", x"00", x"10", x"30", x"20", x"60", x"44", x"84", x"8C", x"81", x"87", x"87", x"87", x"CF", x"CF", x"CF", x"CF", x"00", x"06", x"06", x"06", x"0C", x"0C", x"0C", x"0C", x"F0", x"E0", x"E0", x"E0", x"C1", x"C1", x"C3", x"C3", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"07", x"3F", x"7F", x"FF", x"FF", x"F9", x"F1", x"F0", x"00", x"20", x"40", x"83", x"87", x"01", x"01", x"00", x"C0", x"F0", x"F8", x"FB", x"FB", x"FF", x"FF", x"0F", x"00", x"00", x"00", x"82", x"82", x"FC", x"FC", x"0C", x"1F", x"7F", x"FF", x"FF", x"FF", x"E3", x"C1", x"C1", x"00", x"00", x"00", x"0E", x"1F", x"03", x"01", x"01", 
															x"81", x"C7", x"E7", x"E7", x"F7", x"FF", x"FF", x"FF", x"00", x"06", x"04", x"04", x"04", x"0C", x"08", x"08", x"F0", x"F3", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"00", x"03", x"06", x"06", x"0C", x"0C", x"48", x"48", x"FC", x"FC", x"FC", x"F8", x"F8", x"F8", x"F8", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F8", x"18", x"18", x"18", 
															x"03", x"0F", x"0F", x"0F", x"1F", x"1F", x"1F", x"1F", x"00", x"0C", x"0C", x"0C", x"18", x"18", x"18", x"18", x"FF", x"FB", x"F7", x"07", x"0F", x"1F", x"1F", x"3E", x"01", x"03", x"F6", x"04", x"0C", x"18", x"1F", x"3E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"07", x"0C", x"00", x"00", x"00", x"3E", x"7E", x"07", x"07", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BF", x"BF", x"18", x"18", x"18", x"18", x"10", x"10", x"BF", x"BF", x"83", x"83", x"83", x"FF", x"FD", x"FD", x"F8", x"F8", x"03", x"03", x"03", x"01", x"01", x"01", x"F8", x"F8", x"F0", x"F0", x"F8", x"FF", x"FF", x"FF", x"FF", x"3E", x"00", x"00", x"00", x"80", x"80", x"E0", x"FF", x"3E", x"0F", x"7F", x"FF", x"FF", x"E7", x"C7", x"83", x"00", x"0C", x"0C", x"0C", x"0E", x"06", x"47", x"83", x"00", x"C1", x"C3", x"E7", x"FF", x"FF", x"FF", x"FE", x"F8", x"01", x"02", x"04", x"00", x"00", x"81", x"FE", x"F8", 
															x"FF", x"FF", x"FF", x"DF", x"BF", x"3F", x"79", x"79", x"08", x"18", x"10", x"10", x"31", x"21", x"79", x"79", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E7", x"C7", x"41", x"C1", x"C3", x"C3", x"C2", x"C6", x"E7", x"C7", x"F0", x"F0", x"F0", x"E0", x"E0", x"E0", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"1F", x"FF", x"FF", x"FF", x"FF", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"E0", x"E0", x"C0", x"C0", x"80", 
															x"3F", x"3F", x"3F", x"3F", x"7E", x"7E", x"7C", x"7C", x"30", x"30", x"30", x"30", x"60", x"60", x"7C", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E9", x"4F", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"41", x"32", x"8A", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C7", x"24", x"2F", x"48", x"88", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"BD", x"11", x"11", x"21", x"21", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"29", x"52", x"E7", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"9E", x"92", x"BC", x"A2", x"A2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"40", x"F0", x"80", x"F0", x"00", x"00", 
															x"03", x"0F", x"1F", x"3F", x"3F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"F8", x"FC", x"FC", x"FE", x"FE", x"FE", x"20", x"08", x"04", x"02", x"02", x"01", x"01", x"01", x"7F", x"7F", x"7F", x"3F", x"3F", x"1F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"FE", x"FE", x"FE", x"FC", x"FC", x"F8", x"E0", x"00", x"01", x"01", x"01", x"02", x"02", x"04", x"18", x"E0", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"8F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"1F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"F8", x"F8", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"44", x"C6", x"C6", x"C6", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"2C", x"4C", x"8C", x"FE", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"78", x"C4", x"E4", x"7C", x"9E", x"86", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"38", x"44", x"C6", x"C6", x"C6", x"44", x"38", x"00", x"38", x"44", x"C6", x"C6", x"C6", x"44", x"38", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"E6", x"DA", x"DE", x"DE", x"DE", x"DE", x"DA", x"E6", x"19", x"25", x"21", x"21", x"21", x"21", x"25", x"19", x"D8", x"DB", x"DB", x"18", x"DB", x"DB", x"DB", x"D8", x"27", x"24", x"24", x"E7", x"24", x"24", x"24", x"27", x"66", x"DA", x"DE", x"DE", x"DE", x"DE", x"DA", x"66", x"99", x"25", x"21", x"21", x"21", x"21", x"25", x"99", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"40", x"C0", x"CE", x"C6", x"66", x"3E", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"FE", x"C6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"18", x"18", x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"CC", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"CC", x"D8", x"F0", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"44", x"6C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"D6", x"FE", x"FE", x"6C", x"44", x"00", 
															x"1F", x"07", x"03", x"01", x"01", x"01", x"00", x"00", x"E0", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"24", x"3C", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"08", x"10", x"00", x"DE", x"BE", x"BE", x"7E", x"BE", x"BE", x"DE", x"DE", x"21", x"41", x"41", x"81", x"41", x"41", x"21", x"21", x"39", x"D6", x"D6", x"D6", x"36", x"F6", x"F6", x"F9", x"C6", x"29", x"29", x"29", x"C9", x"09", x"09", x"06", x"8B", x"D9", x"D9", x"DA", x"DA", x"DB", x"DB", x"8B", x"74", x"26", x"26", x"25", x"25", x"24", x"24", x"74", x"43", x"6F", x"6F", x"6F", x"6F", x"6F", x"6F", x"6F", x"BC", x"90", x"90", x"90", x"90", x"90", x"90", x"90", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"FF", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"03", x"02", x"13", x"0A", x"05", x"04", x"00", x"00", x"01", x"00", x"11", x"0D", x"06", x"0B", x"00", x"00", x"40", x"00", x"C0", x"30", x"60", x"A0", x"00", x"40", x"40", x"00", x"80", x"A0", x"C0", x"D0", x"01", x"83", x"62", x"3F", x"15", x"1A", x"3D", x"E2", x"01", x"8B", x"63", x"3F", x"1F", x"1D", x"3F", x"F5", x"00", x"06", x"40", x"98", x"30", x"E0", x"70", x"A0", x"00", x"06", x"64", x"9C", x"90", x"F0", x"F0", x"F4", x"00", x"08", x"00", x"28", x"10", x"05", x"2C", x"09", x"00", x"0C", x"03", x"3A", x"15", x"15", x"2E", x"0D", x"08", x"10", x"00", x"A0", x"24", x"40", x"A8", x"00", x"8C", x"50", x"A8", x"B0", x"64", x"D2", x"E8", x"90", x"0F", x"17", x"1F", x"1F", x"1F", x"1F", x"19", x"13", x"0F", x"1F", x"0F", x"0F", x"0F", x"1F", x"1E", x"1C", x"C0", x"60", x"E0", x"E0", x"F0", x"F0", x"F0", x"F8", x"80", x"C0", x"80", x"80", x"80", x"C0", x"C0", x"40", 
															x"00", x"00", x"00", x"00", x"01", x"07", x"06", x"02", x"00", x"01", x"03", x"07", x"06", x"00", x"01", x"01", x"00", x"00", x"10", x"08", x"80", x"C0", x"D8", x"18", x"00", x"80", x"E0", x"D0", x"70", x"30", x"30", x"E8", x"00", x"00", x"00", x"08", x"0F", x"0F", x"0F", x"0C", x"07", x"0F", x"1F", x"1F", x"18", x"18", x"10", x"17", x"40", x"30", x"18", x"18", x"98", x"D8", x"DC", x"5E", x"80", x"C0", x"E0", x"E0", x"60", x"20", x"20", x"A0", x"00", x"10", x"30", x"10", x"10", x"16", x"2F", x"0F", x"00", x"0F", x"1F", x"3F", x"3F", x"30", x"10", x"10", x"80", x"C0", x"60", x"30", x"30", x"30", x"78", x"78", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"80", x"80", x"07", x"00", x"18", x"00", x"1F", x"1F", x"1C", x"18", x"00", x"0F", x"07", x"1F", x"10", x"18", x"07", x"07", x"E0", x"70", x"B0", x"30", x"B0", x"78", x"FC", x"FC", x"00", x"80", x"40", x"C0", x"40", x"80", x"00", x"00", 
															x"1A", x"07", x"0D", x"24", x"00", x"04", x"00", x"00", x"1D", x"06", x"0B", x"24", x"00", x"04", x"00", x"00", x"74", x"68", x"D0", x"C0", x"40", x"00", x"00", x"00", x"B4", x"E0", x"90", x"C0", x"00", x"00", x"00", x"00", x"07", x"0F", x"0D", x"14", x"28", x"20", x"00", x"00", x"07", x"0F", x"0F", x"1C", x"38", x"20", x"40", x"00", x"3C", x"A0", x"60", x"D0", x"B0", x"98", x"80", x"02", x"7C", x"A0", x"E0", x"F0", x"B0", x"D8", x"84", x"02", x"02", x"05", x"20", x"01", x"00", x"02", x"00", x"04", x"0B", x"07", x"28", x"01", x"01", x"02", x"00", x"04", x"40", x"C0", x"20", x"00", x"10", x"08", x"00", x"00", x"C8", x"E0", x"60", x"00", x"10", x"08", x"00", x"00", x"17", x"17", x"17", x"17", x"1F", x"1F", x"1F", x"1F", x"18", x"1F", x"1F", x"1F", x"0F", x"08", x"0F", x"1F", x"F8", x"F8", x"F8", x"F8", x"F8", x"F0", x"F0", x"F0", x"40", x"40", x"40", x"40", x"80", x"80", x"80", x"C0", 
															x"06", x"00", x"01", x"03", x"03", x"03", x"03", x"00", x"01", x"07", x"07", x"07", x"06", x"06", x"04", x"00", x"F0", x"50", x"18", x"C0", x"90", x"20", x"D4", x"00", x"50", x"F0", x"E8", x"30", x"68", x"D8", x"24", x"00", x"0C", x"0C", x"0F", x"07", x"00", x"0C", x"00", x"0F", x"17", x"1B", x"10", x"18", x"1F", x"13", x"1F", x"10", x"5E", x"5E", x"DE", x"9C", x"18", x"D8", x"18", x"DC", x"A0", x"A0", x"20", x"60", x"E0", x"20", x"E0", x"20", x"08", x"08", x"28", x"3F", x"1F", x"1F", x"10", x"1F", x"1F", x"1F", x"1F", x"30", x"30", x"30", x"2F", x"20", x"7C", x"7C", x"7C", x"7C", x"38", x"38", x"30", x"B8", x"80", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"40", x"18", x"00", x"00", x"1F", x"07", x"00", x"00", x"0F", x"07", x"1F", x"1F", x"00", x"18", x"1F", x"0F", x"00", x"FC", x"3C", x"3C", x"F8", x"B8", x"30", x"70", x"F0", x"00", x"C0", x"C0", x"00", x"40", x"C0", x"80", x"00", 
															x"00", x"1F", x"2F", x"2F", x"2F", x"27", x"3F", x"1F", x"00", x"0F", x"1F", x"3F", x"3F", x"30", x"10", x"10", x"00", x"00", x"20", x"30", x"30", x"30", x"18", x"18", x"00", x"00", x"E0", x"D0", x"D0", x"D0", x"F8", x"F8", x"08", x"08", x"10", x"10", x"10", x"1E", x"0F", x"11", x"1F", x"3F", x"3F", x"3F", x"3F", x"31", x"20", x"2E", x"C0", x"60", x"60", x"60", x"70", x"70", x"70", x"78", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"0F", x"1F", x"1F", x"2F", x"2F", x"2F", x"3F", x"1F", x"0F", x"1F", x"1F", x"3F", x"3D", x"38", x"30", x"17", x"80", x"40", x"00", x"20", x"30", x"30", x"38", x"78", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"00", x"00", x"00", x"00", x"01", x"0E", x"15", x"2F", x"00", x"00", x"00", x"00", x"01", x"0F", x"1F", x"39", x"38", x"DC", x"BC", x"7E", x"FE", x"FE", x"FE", x"FC", x"38", x"FC", x"FC", x"FE", x"3E", x"1E", x"8C", x"D0", 
															x"00", x"00", x"00", x"00", x"03", x"0E", x"1B", x"37", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"39", x"00", x"00", x"0E", x"27", x"5F", x"FF", x"FF", x"FF", x"00", x"00", x"0E", x"3F", x"7F", x"DF", x"8F", x"CF", x"00", x"00", x"00", x"F8", x"FF", x"E7", x"F8", x"FF", x"00", x"00", x"00", x"F8", x"FF", x"7F", x"77", x"73", x"00", x"00", x"00", x"F0", x"F8", x"FE", x"BE", x"FE", x"00", x"00", x"00", x"60", x"F0", x"F8", x"7C", x"3C", x"7C", x"FE", x"FF", x"7F", x"BF", x"FF", x"77", x"3F", x"7C", x"FE", x"FE", x"FB", x"F1", x"E3", x"6F", x"3E", x"00", x"00", x"00", x"C0", x"E0", x"38", x"98", x"CC", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"70", x"00", x"18", x"7E", x"7E", x"FF", x"FF", x"FF", x"BF", x"00", x"18", x"7E", x"7E", x"F9", x"F1", x"F3", x"E3", x"00", x"00", x"00", x"F0", x"FC", x"06", x"43", x"E1", x"00", x"00", x"00", x"00", x"00", x"F8", x"FC", x"3E", 
															x"17", x"17", x"37", x"0F", x"2F", x"2F", x"3F", x"3F", x"1F", x"1F", x"1F", x"30", x"30", x"30", x"2F", x"10", x"7C", x"7C", x"7C", x"3C", x"38", x"78", x"F0", x"60", x"FC", x"FC", x"FC", x"DC", x"D8", x"D8", x"50", x"A0", x"11", x"11", x"11", x"0E", x"1F", x"00", x"00", x"1F", x"2E", x"2E", x"2E", x"31", x"20", x"3F", x"3F", x"20", x"78", x"78", x"78", x"78", x"70", x"60", x"60", x"60", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"1B", x"1B", x"1F", x"37", x"3F", x"3F", x"3F", x"3F", x"17", x"17", x"10", x"38", x"2F", x"2F", x"3F", x"20", x"78", x"78", x"78", x"30", x"B0", x"B0", x"38", x"D0", x"80", x"80", x"80", x"C0", x"40", x"40", x"C0", x"20", x"7F", x"7F", x"7F", x"1F", x"0F", x"0F", x"07", x"03", x"78", x"7C", x"1E", x"0F", x"07", x"07", x"03", x"03", x"98", x"38", x"10", x"30", x"30", x"60", x"C0", x"80", x"E0", x"C0", x"E0", x"C0", x"C0", x"80", x"00", x"00", 
															x"7F", x"7F", x"3F", x"1F", x"0F", x"0F", x"0F", x"0F", x"3C", x"3C", x"0E", x"0E", x"07", x"07", x"07", x"06", x"FD", x"F7", x"CF", x"DE", x"F8", x"B0", x"60", x"C0", x"CE", x"78", x"70", x"60", x"C0", x"C0", x"80", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"F8", x"00", x"00", x"73", x"73", x"77", x"FF", x"F8", x"00", x"00", x"00", x"FE", x"FE", x"FC", x"F8", x"F0", x"60", x"00", x"00", x"3C", x"3C", x"78", x"F0", x"60", x"00", x"00", x"00", x"17", x"1B", x"1F", x"1F", x"0F", x"07", x"07", x"03", x"1C", x"1C", x"19", x"1F", x"0F", x"07", x"06", x"02", x"FC", x"FC", x"F8", x"E0", x"C0", x"80", x"80", x"00", x"78", x"F8", x"E0", x"C0", x"80", x"00", x"00", x"00", x"5B", x"1F", x"07", x"02", x"03", x"01", x"00", x"00", x"7E", x"1E", x"06", x"03", x"03", x"01", x"00", x"00", x"FF", x"FC", x"F8", x"78", x"B0", x"F8", x"78", x"70", x"78", x"78", x"F0", x"F0", x"E0", x"F0", x"70", x"00", 
															x"00", x"00", x"00", x"1F", x"3F", x"7F", x"FF", x"FF", x"00", x"00", x"00", x"18", x"3F", x"7F", x"F3", x"F3", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"7C", x"FC", x"B8", x"38", x"38", x"00", x"10", x"00", x"00", x"1F", x"10", x"10", x"10", x"1F", x"1F", x"3F", x"3F", x"20", x"2F", x"3F", x"3F", x"70", x"78", x"38", x"38", x"BE", x"BE", x"3E", x"3E", x"80", x"80", x"C0", x"C0", x"40", x"40", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"D5", x"D5", x"D5", x"D5", x"D5", x"D5", x"81", x"42", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"E0", x"C0", x"78", x"78", x"78", x"78", x"78", x"78", x"60", x"C0", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"04", x"1C", x"1C", x"1C", x"1E", x"3E", x"7E", x"00", x"18", x"18", x"18", x"18", x"1C", x"0C", x"04", x"03", x"07", x"04", x"08", x"08", x"0C", x"07", x"03", x"00", x"03", x"07", x"0B", x"03", x"07", x"03", x"00", x"C0", x"E0", x"20", x"50", x"10", x"30", x"E0", x"C0", x"00", x"C0", x"E0", x"F0", x"E0", x"E0", x"C0", x"00", x"3F", x"3F", x"3F", x"3F", x"3F", x"20", x"2F", x"32", x"24", x"25", x"25", x"25", x"24", x"20", x"20", x"2D", x"F8", x"FC", x"FE", x"FF", x"FF", x"3F", x"9F", x"CF", x"80", x"48", x"54", x"54", x"94", x"08", x"00", x"00", x"12", x"14", x"7C", x"7C", x"7C", x"7C", x"7C", x"3C", x"6C", x"68", x"00", x"68", x"68", x"68", x"68", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"38", x"30", x"00", x"40", x"00", x"00", x"00", 
															x"FF", x"EC", x"FF", x"7F", x"3F", x"18", x"00", x"00", x"F3", x"FB", x"7F", x"3F", x"18", x"00", x"00", x"00", x"FE", x"7E", x"DE", x"FE", x"7E", x"00", x"00", x"00", x"38", x"B8", x"F8", x"7C", x"3C", x"00", x"00", x"00", x"16", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"09", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"EC", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"55", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D5", x"D5", x"D5", x"D5", x"D5", x"D5", x"81", x"81", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"E0", x"C0", x"78", x"78", x"78", x"78", x"78", x"78", x"60", x"40", 
															x"00", x"03", x"03", x"03", x"03", x"01", x"00", x"00", x"03", x"03", x"03", x"03", x"01", x"00", x"00", x"00", x"7E", x"7A", x"02", x"43", x"A5", x"29", x"32", x"2A", x"00", x"04", x"3C", x"3C", x"7E", x"FE", x"FF", x"FF", x"26", x"01", x"01", x"02", x"02", x"06", x"C6", x"3E", x"FD", x"FE", x"FE", x"FC", x"FC", x"F8", x"3C", x"2C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"03", x"03", x"1F", x"3F", x"3F", x"3F", x"3F", x"1F", x"1F", x"07", x"08", x"0D", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"F8", x"FC", x"FC", x"FC", x"F8", x"F0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"0F", x"06", x"03", x"01", x"00", x"00", x"01", x"02", x"06", x"02", x"01", x"00", x"00", x"EC", x"FE", x"BC", x"F8", x"F0", x"E0", x"C0", x"00", x"A0", x"98", x"80", x"60", x"00", x"80", x"00", x"00", 
															x"00", x"1F", x"1F", x"13", x"1F", x"1F", x"1F", x"1F", x"00", x"00", x"0D", x"01", x"0D", x"0D", x"0D", x"00", x"00", x"F8", x"F8", x"48", x"F8", x"F8", x"F8", x"F8", x"00", x"00", x"B0", x"00", x"B0", x"B0", x"B0", x"00", x"01", x"3F", x"3F", x"03", x"3F", x"3F", x"01", x"FF", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"39", x"11", x"01", x"01", x"29", x"39", x"39", x"FF", x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"03", x"39", x"39", x"39", x"03", x"3F", x"3F", x"FF", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"81", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"FF", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"07", x"0F", x"0F", x"0F", x"0F", x"07", x"00", x"07", x"0F", x"1F", x"1F", x"1F", x"1C", x"08", x"00", x"20", x"D0", x"E8", x"E8", x"E8", x"E8", x"D0", x"00", x"C0", x"E0", x"F0", x"F0", x"F0", x"70", x"20", 
															x"03", x"0F", x"1F", x"1B", x"17", x"17", x"2F", x"2F", x"00", x"00", x"00", x"04", x"08", x"08", x"10", x"10", x"E0", x"F0", x"F8", x"F8", x"FC", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"33", x"33", x"CF", x"CF", x"33", x"32", x"CE", x"CE", x"CC", x"CC", x"30", x"30", x"CC", x"CD", x"31", x"31", x"33", x"33", x"FF", x"FF", x"07", x"7B", x"7F", x"7F", x"CC", x"CC", x"00", x"00", x"F8", x"84", x"80", x"80", x"33", x"33", x"FF", x"FF", x"83", x"39", x"39", x"39", x"CC", x"CC", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"33", x"33", x"FF", x"FF", x"F7", x"EB", x"DD", x"DD", x"CC", x"CC", x"00", x"00", x"08", x"14", x"22", x"22", x"33", x"33", x"FF", x"FF", x"CF", x"CF", x"CF", x"CF", x"CC", x"CC", x"00", x"00", x"30", x"30", x"30", x"30", x"33", x"33", x"CC", x"CC", x"F3", x"F3", x"CC", x"CC", x"CC", x"CC", x"33", x"33", x"0C", x"0C", x"33", x"33", 
															x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FE", x"FC", x"F8", x"E0", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"99", x"99", x"DB", x"C3", x"E7", x"E7", x"E7", x"FF", x"66", x"66", x"24", x"3C", x"18", x"18", x"18", x"00", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"0C", x"0C", x"08", x"0F", x"17", x"10", x"10", x"1F", x"0B", x"0B", x"0F", x"08", x"18", x"1F", x"1F", x"1F", x"7C", x"7C", x"3C", x"FC", x"DC", x"1C", x"1C", x"F8", x"A0", x"A0", x"E0", x"20", x"30", x"F0", x"F0", x"F0", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"A7", x"EF", x"CA", x"EA", x"AA", x"AA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"14", x"17", x"A7", x"A5", x"C5", x"C5", x"85", x"32", x"32", x"CE", x"CF", x"33", x"33", x"CC", x"CC", x"CD", x"CD", x"31", x"30", x"CC", x"CC", x"33", x"33", x"43", x"73", x"73", x"07", x"FF", x"FF", x"CC", x"CC", x"BC", x"8C", x"8C", x"F8", x"00", x"00", x"33", x"33", x"39", x"39", x"39", x"83", x"FF", x"FF", x"CC", x"CC", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"33", x"33", x"80", x"9C", x"9C", x"9C", x"FF", x"FF", x"CC", x"CC", x"7F", x"63", x"63", x"63", x"00", x"00", x"33", x"33", x"CF", x"CF", x"CF", x"C0", x"FF", x"FF", x"CC", x"CC", x"30", x"30", x"30", x"3F", x"00", x"00", x"33", x"33", x"F3", x"F3", x"CC", x"4C", x"F3", x"F3", x"CC", x"CC", x"0C", x"0C", x"33", x"B3", x"0C", x"0C", x"33", x"33", 
															x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"7E", x"3C", x"00", x"3C", x"7E", x"FF", x"E7", x"C3", x"C3", x"7E", x"FF", x"87", x"BB", x"BA", x"BA", x"86", x"BE", x"BE", x"00", x"78", x"44", x"45", x"45", x"79", x"41", x"41", x"FF", x"BB", x"5B", x"EB", x"0B", x"EB", x"EB", x"EC", x"00", x"44", x"A4", x"14", x"F4", x"14", x"14", x"13", x"FF", x"B1", x"AE", x"AF", x"A1", x"BE", x"AE", x"71", x"00", x"4E", x"51", x"50", x"5E", x"41", x"51", x"8E", x"FF", x"83", x"BF", x"BF", x"87", x"BF", x"BF", x"83", x"00", x"7C", x"40", x"40", x"78", x"40", x"40", x"7C", x"00", x"00", x"10", x"10", x"10", x"00", x"07", x"0F", x"0F", x"1F", x"0F", x"0F", x"0F", x"1F", x"1E", x"1C", x"60", x"30", x"70", x"70", x"70", x"38", x"3C", x"B0", x"80", x"C0", x"80", x"80", x"80", x"C0", x"C0", x"40", x"4A", x"6A", x"5A", x"4A", x"4A", x"00", x"0F", x"12", x"4A", x"6A", x"5A", x"4A", x"4A", x"00", x"00", x"0D", 
															x"67", x"94", x"87", x"94", x"67", x"00", x"80", x"C0", x"67", x"94", x"87", x"94", x"67", x"00", x"00", x"00", x"B2", x"18", x"C7", x"EF", x"4F", x"5F", x"9F", x"1F", x"00", x"00", x"00", x"02", x"04", x"06", x"00", x"00", x"13", x"27", x"CE", x"E0", x"F3", x"F3", x"F8", x"F8", x"00", x"00", x"00", x"80", x"40", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"F8", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"17", x"03", x"00", x"00", x"07", x"07", x"08", x"0F", x"08", x"1C", x"1F", x"1F", x"18", x"18", x"17", x"10", x"B8", x"18", x"18", x"18", x"9C", x"9C", x"5C", x"C0", x"40", x"E0", x"E0", x"E0", x"60", x"60", x"A0", 
															x"3C", x"3C", x"3C", x"7E", x"7E", x"7E", x"00", x"00", x"7E", x"7E", x"42", x"C3", x"FF", x"FF", x"FF", x"81", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"80", x"9F", x"90", x"9E", x"90", x"90", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"22", x"22", x"22", x"22", x"1C", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"7C", x"40", x"7C", x"40", x"7C", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"01", x"81", x"81", x"81", x"81", x"F9", x"FF", x"0F", x"0F", x"0F", x"18", x"13", x"10", x"00", x"0F", x"1C", x"18", x"18", x"0F", x"0C", x"0F", x"1F", x"10", x"B0", x"B0", x"B0", x"78", x"78", x"78", x"38", x"B8", x"40", x"40", x"40", x"80", x"80", x"80", x"C0", x"40", x"1F", x"3F", x"3F", x"3F", x"3F", x"1F", x"1F", x"07", x"08", x"0D", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"E0", x"F0", x"F8", x"FC", x"FC", x"FC", x"F8", x"F0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"3F", x"3F", x"3F", x"1F", x"19", x"33", x"26", x"1F", x"00", x"00", x"00", x"00", x"E6", x"4C", x"19", x"00", x"FC", x"FC", x"F8", x"E8", x"98", x"30", x"67", x"FE", x"00", x"00", x"00", x"00", x"66", x"CC", x"98", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"0B", x"0B", x"0C", x"0F", x"07", x"00", x"00", x"08", x"17", x"17", x"13", x"10", x"18", x"1F", x"1F", x"0F", x"5E", x"5C", x"DC", x"D8", x"98", x"18", x"10", x"70", x"A0", x"A0", x"20", x"20", x"60", x"E0", x"E0", x"C0");
	
	constant PINBALL_CHR_ROM : CHR_ROM_ARRAY := (x"00", x"00", x"00", x"07", x"05", x"05", x"0F", x"07", x"00", x"07", x"0F", x"07", x"07", x"07", x"0F", x"07", x"00", x"00", x"00", x"80", x"80", x"80", x"40", x"C0", x"00", x"C0", x"E0", x"E0", x"E0", x"E0", x"F6", x"FC", x"03", x"21", x"63", x"7F", x"1F", x"04", x"03", x"03", x"03", x"21", x"61", x"60", x"00", x"03", x"00", x"00", x"80", x"C0", x"E0", x"E0", x"B0", x"3C", x"DC", x"D0", x"F8", x"3C", x"10", x"08", x"00", x"8C", x"1C", x"10", x"07", x"07", x"0F", x"0F", x"0F", x"1F", x"00", x"00", x"00", x"00", x"00", x"01", x"0E", x"00", x"0C", x"1C", x"E0", x"F8", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"00", x"10", x"60", x"8C", x"1C", x"08", x"08", x"00", x"00", x"00", x"07", x"05", x"05", x"0F", x"07", x"03", x"07", x"0F", x"07", x"07", x"07", x"0F", x"07", x"03", x"00", x"00", x"80", x"80", x"80", x"40", x"C0", x"80", x"C0", x"E0", x"E0", x"E0", x"E0", x"F0", x"F8", x"FC", 
															x"01", x"03", x"07", x"07", x"0C", x"07", x"03", x"07", x"01", x"01", x"00", x"00", x"0F", x"04", x"00", x"00", x"C0", x"E0", x"E0", x"F0", x"70", x"E0", x"C0", x"C0", x"34", x"10", x"18", x"04", x"80", x"C0", x"C0", x"80", x"07", x"0F", x"0F", x"0F", x"1F", x"01", x"00", x"00", x"00", x"00", x"00", x"0F", x"00", x"06", x"0E", x"01", x"E0", x"E0", x"F0", x"F0", x"F8", x"E0", x"00", x"00", x"00", x"00", x"00", x"70", x"C0", x"00", x"C0", x"C0", x"01", x"01", x"03", x"12", x"3D", x"3F", x"07", x"03", x"01", x"00", x"00", x"11", x"32", x"30", x"00", x"00", x"C0", x"E0", x"E0", x"E0", x"C0", x"F0", x"30", x"C0", x"30", x"18", x"0C", x"00", x"20", x"30", x"F0", x"00", x"07", x"2F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"08", x"06", x"11", x"78", x"18", x"00", x"00", x"E0", x"E0", x"E0", x"F8", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"90", x"60", x"18", x"30", x"60", 
															x"01", x"03", x"07", x"07", x"0C", x"3B", x"0B", x"07", x"01", x"01", x"00", x"00", x"03", x"38", x"08", x"00", x"C0", x"E0", x"F0", x"F8", x"38", x"DE", x"CE", x"E8", x"30", x"18", x"04", x"00", x"80", x"0E", x"0E", x"08", x"07", x"0F", x"0F", x"0F", x"1F", x"07", x"00", x"00", x"00", x"00", x"00", x"0C", x"03", x"00", x"06", x"0E", x"E0", x"E0", x"F0", x"F0", x"F8", x"F0", x"00", x"00", x"00", x"00", x"00", x"10", x"E0", x"00", x"60", x"70", x"00", x"00", x"00", x"0E", x"0B", x"1B", x"3F", x"31", x"28", x"3F", x"1F", x"0F", x"0F", x"1F", x"3F", x"31", x"00", x"00", x"00", x"00", x"00", x"40", x"C0", x"80", x"00", x"80", x"C0", x"C0", x"C0", x"EC", x"F8", x"F0", x"19", x"0F", x"1F", x"3F", x"F7", x"E7", x"20", x"03", x"19", x"0F", x"02", x"00", x"C0", x"E0", x"23", x"00", x"E0", x"FE", x"FF", x"CC", x"C4", x"B0", x"78", x"FE", x"98", x"06", x"07", x"04", x"04", x"40", x"80", x"04", 
															x"07", x"07", x"07", x"0F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"FC", x"FC", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"08", x"10", x"66", x"87", x"23", x"60", x"20", x"00", x"00", x"00", x"00", x"00", x"07", x"05", x"05", x"0F", x"00", x"02", x"07", x"17", x"1F", x"0F", x"07", x"0F", x"00", x"00", x"00", x"00", x"C0", x"60", x"50", x"F0", x"80", x"80", x"E0", x"F0", x"F2", x"F4", x"FE", x"FC", x"0C", x"0C", x"0E", x"0F", x"07", x"26", x"3A", x"3F", x"0F", x"0F", x"07", x"01", x"00", x"01", x"01", x"01", x"60", x"70", x"78", x"F8", x"F0", x"E6", x"DE", x"FE", x"FC", x"E8", x"E0", x"C0", x"00", x"00", x"24", x"C4", x"1F", x"0F", x"07", x"0F", x"0E", x"0C", x"00", x"00", x"03", x"01", x"00", x"1F", x"1E", x"1C", x"18", x"00", x"FC", x"F8", x"F0", x"78", x"78", x"30", x"00", x"00", x"88", x"00", x"16", x"7E", x"7E", x"32", x"00", x"00", 
															x"00", x"00", x"07", x"0D", x"07", x"03", x"07", x"1F", x"00", x"0F", x"07", x"0F", x"07", x"03", x"01", x"00", x"00", x"00", x"C0", x"A0", x"E0", x"C0", x"F0", x"F8", x"00", x"F0", x"F0", x"FA", x"FC", x"F8", x"8C", x"06", x"7F", x"10", x"07", x"0F", x"1F", x"1F", x"1F", x"00", x"70", x"13", x"00", x"00", x"00", x"1F", x"00", x"3C", x"DC", x"0E", x"EC", x"F0", x"F8", x"F8", x"F8", x"00", x"00", x"CE", x"0C", x"00", x"00", x"F8", x"00", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"09", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"99", x"FF", x"00", x"01", x"01", x"00", x"07", x"00", x"00", x"00", x"00", x"07", x"07", x"1F", x"07", x"FF", x"99", x"FF", x"E0", x"E0", x"C0", x"C0", x"00", x"00", x"00", x"60", x"E0", x"E0", x"C0", x"20", x"E0", 
															x"3A", x"7E", x"3E", x"1E", x"0E", x"02", x"02", x"02", x"01", x"09", x"3D", x"01", x"01", x"07", x"0F", x"1F", x"30", x"30", x"38", x"30", x"00", x"00", x"00", x"00", x"D0", x"D0", x"F8", x"D0", x"C0", x"E0", x"E0", x"E0", x"06", x"07", x"1F", x"1F", x"0F", x"0F", x"00", x"00", x"1F", x"1F", x"1B", x"1F", x"0F", x"0F", x"07", x"0F", x"20", x"20", x"E0", x"F0", x"F8", x"78", x"00", x"00", x"E0", x"E0", x"E8", x"FC", x"FE", x"7A", x"00", x"00", x"FF", x"99", x"FF", x"00", x"00", x"00", x"03", x"1D", x"00", x"00", x"00", x"03", x"03", x"0F", x"03", x"1D", x"FF", x"99", x"FF", x"F0", x"E0", x"60", x"80", x"10", x"00", x"00", x"70", x"F0", x"E0", x"90", x"F0", x"F0", x"3F", x"1F", x"0F", x"07", x"01", x"01", x"01", x"03", x"04", x"1E", x"00", x"00", x"03", x"07", x"0F", x"0F", x"18", x"1C", x"18", x"00", x"00", x"00", x"80", x"80", x"E8", x"FC", x"E8", x"E0", x"F0", x"F0", x"F0", x"F0", 
															x"0F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"00", x"0D", x"0F", x"0B", x"07", x"07", x"0F", x"00", x"00", x"90", x"F0", x"F0", x"F0", x"F0", x"E0", x"00", x"00", x"F0", x"F0", x"F0", x"F0", x"F0", x"E0", x"E0", x"E0", x"3F", x"1F", x"0F", x"07", x"00", x"00", x"00", x"01", x"04", x"1E", x"00", x"00", x"01", x"03", x"07", x"07", x"18", x"1C", x"18", x"00", x"80", x"80", x"80", x"88", x"E8", x"FC", x"E8", x"F0", x"F0", x"F0", x"F0", x"F8", x"07", x"07", x"0F", x"0F", x"07", x"00", x"00", x"00", x"06", x"07", x"2F", x"3F", x"1F", x"08", x"00", x"00", x"D8", x"F8", x"F8", x"FC", x"FC", x"38", x"00", x"00", x"F8", x"F8", x"F8", x"FC", x"FE", x"3E", x"06", x"0C", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"7F", x"00", x"7F", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", 
															x"00", x"00", x"00", x"00", x"00", x"3C", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"3C", x"00", x"3C", x"00", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"3F", x"40", x"40", x"40", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"0E", x"1C", x"18", x"10", x"03", x"0F", x"1F", x"39", x"71", x"63", x"E7", x"EF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"F8", x"FC", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C3", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"81", x"C3", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"7F", x"7F", x"3F", x"1F", x"0F", x"03", 
															x"02", x"02", x"03", x"03", x"03", x"03", x"02", x"02", x"02", x"02", x"03", x"03", x"03", x"03", x"02", x"02", x"02", x"06", x"04", x"0C", x"0C", x"08", x"08", x"00", x"0E", x"06", x"04", x"0C", x"0C", x"08", x"08", x"00", x"04", x"04", x"0C", x"08", x"08", x"00", x"00", x"00", x"0C", x"04", x"0C", x"08", x"08", x"00", x"00", x"00", x"06", x"06", x"03", x"03", x"03", x"03", x"06", x"06", x"06", x"06", x"03", x"0F", x"0F", x"03", x"06", x"06", x"06", x"06", x"0C", x"0C", x"0C", x"08", x"08", x"08", x"06", x"06", x"0C", x"0C", x"0C", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"38", x"1E", x"0F", x"00", x"00", x"00", x"00", x"00", x"38", x"1E", x"0F", x"38", x"18", x"0C", x"0C", x"06", x"02", x"00", x"00", x"38", x"38", x"0C", x"0C", x"06", x"02", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"03", x"03", x"00", x"00", x"01", x"01", x"03", x"03", x"03", x"03", 
															x"03", x"06", x"06", x"0E", x"1C", x"38", x"70", x"40", x"03", x"0E", x"0E", x"0E", x"1C", x"38", x"70", x"40", x"00", x"40", x"20", x"30", x"18", x"1C", x"0E", x"07", x"00", x"40", x"20", x"30", x"18", x"1C", x"0E", x"07", x"38", x"1C", x"0C", x"0C", x"06", x"06", x"06", x"06", x"38", x"1C", x"1C", x"3C", x"16", x"06", x"06", x"06", x"03", x"03", x"03", x"03", x"01", x"01", x"00", x"00", x"03", x"03", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"00", x"10", x"08", x"08", x"0C", x"06", x"06", x"00", x"00", x"10", x"08", x"08", x"0C", x"06", x"06", x"30", x"38", x"18", x"0C", x"0C", x"0C", x"0C", x"0C", x"30", x"38", x"18", x"3C", x"1C", x"0C", x"0C", x"0C", x"06", x"06", x"06", x"06", x"06", x"02", x"02", x"02", x"06", x"06", x"06", x"06", x"06", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FC", x"F8", x"F0", x"C0", 
															x"00", x"00", x"0C", x"1C", x"14", x"1F", x"3E", x"0E", x"00", x"0F", x"03", x"03", x"03", x"07", x"3F", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"E0", x"E0", x"F8", x"FC", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"1F", x"00", x"00", x"00", x"80", x"C8", x"F8", x"D0", x"30", x"00", x"E0", x"F0", x"78", x"38", x"18", x"10", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"0F", x"1F", x"1F", x"3F", x"3F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"3F", x"1F", x"1F", x"0F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", 
															x"18", x"3C", x"3C", x"3C", x"18", x"00", x"00", x"00", x"18", x"3C", x"3C", x"3C", x"18", x"00", x"00", x"00", x"7B", x"73", x"73", x"73", x"74", x"78", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"00", x"00", x"0F", x"0F", x"00", x"00", x"0F", x"0F", x"00", x"00", x"0F", x"0F", x"00", x"00", x"FE", x"FE", x"00", x"00", x"FE", x"FE", x"00", x"00", x"FE", x"FE", x"00", x"00", x"FE", x"FE", x"00", x"FF", x"FD", x"FD", x"FD", x"F9", x"FB", x"76", x"3C", x"00", x"02", x"02", x"02", x"06", x"04", x"08", x"00", x"10", x"22", x"00", x"00", x"87", x"C6", x"62", x"30", x"00", x"10", x"00", x"86", x"48", x"20", x"18", x"00", x"00", x"03", x"07", x"00", x"00", x"1F", x"1F", x"00", x"00", x"03", x"07", x"00", x"00", x"1F", x"1F", x"00", x"00", x"E0", x"F0", x"80", x"80", x"FC", x"FC", x"00", x"00", x"E0", x"F0", x"00", x"00", x"FC", x"FC", x"00", 
															x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"66", x"C0", x"C0", x"C0", x"66", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"CC", x"C6", x"C6", x"C6", x"CC", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"C6", x"EE", x"FE", x"FE", x"D6", x"C6", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"99", x"A1", x"A1", x"99", x"42", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"60", x"61", x"63", x"67", x"63", x"61", x"60", x"00", x"60", x"61", x"63", x"67", x"63", x"61", x"60", x"00", x"FF", x"EF", x"CF", x"EF", x"EF", x"EF", x"FF", x"00", x"FF", x"EF", x"CF", x"EF", x"EF", x"EF", x"FF", x"00", x"FF", x"C7", x"F7", x"C7", x"DF", x"C7", x"FF", x"00", x"FF", x"C7", x"F7", x"C7", x"DF", x"C7", x"FF", x"00", x"FF", x"C7", x"F7", x"E7", x"F7", x"C7", x"FF", x"00", x"FF", x"C7", x"F7", x"E7", x"F7", x"C7", x"FF", x"00", x"FF", x"F7", x"E7", x"D7", x"C3", x"F7", x"FF", x"00", x"FF", x"F7", x"E7", x"D7", x"C3", x"F7", x"FF", x"00", x"FF", x"C7", x"DF", x"C7", x"F7", x"C7", x"FF", x"00", x"FF", x"C7", x"DF", x"C7", x"F7", x"C7", x"FF", x"00", x"FF", x"C7", x"DF", x"C7", x"D7", x"C7", x"FF", x"00", x"FF", x"C7", x"DF", x"C7", x"D7", x"C7", x"FF", x"00", x"FF", x"C7", x"F7", x"EF", x"EF", x"EF", x"FF", x"00", x"FF", x"C7", x"F7", x"EF", x"EF", x"EF", x"FF", x"00", 
															x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C6", x"C6", x"C6", x"EE", x"7C", x"38", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"60", x"E0", x"E0", x"1C", x"1E", x"1D", x"39", x"3F", x"1F", x"1F", x"1E", x"1C", x"1C", x"1C", x"1C", x"0C", x"04", x"00", x"00", x"03", x"03", x"03", x"23", x"73", x"F3", x"03", x"01", x"00", x"00", x"00", x"00", x"40", x"60", x"00", x"00", x"E0", x"E4", x"F4", x"FF", x"BE", x"98", x"C0", x"E0", 
															x"7F", x"7F", x"78", x"74", x"73", x"73", x"73", x"77", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"78", x"7C", x"7F", x"7F", x"7F", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"1E", x"2E", x"CE", x"CE", x"CE", x"2E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5E", x"CE", x"CE", x"CE", x"2E", x"1E", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"7F", x"7F", x"7F", x"7C", x"78", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DE", x"CE", x"CE", x"CE", x"EE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"56", x"56", x"00", x"00", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"0C", x"18", x"3C", x"7E", x"7E", x"3C", x"00", x"7E", x"FC", x"18", x"3C", x"7E", x"7E", x"3C", x"66", 
															x"00", x"00", x"06", x"06", x"60", x"60", x"70", x"F0", x"0C", x"1E", x"3A", x"78", x"1E", x"1E", x"0E", x"0E", x"38", x"38", x"38", x"1C", x"1C", x"0E", x"00", x"00", x"07", x"07", x"07", x"23", x"63", x"F1", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"00", x"00", x"C0", x"C0", x"E4", x"FE", x"FB", x"C0", x"E0", x"F0", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"04", x"00", x"00", x"00", x"07", x"0F", x"09", x"19", x"1B", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"04", x"00", x"00", x"00", x"07", x"0F", x"09", x"19", x"1B", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"1F", x"0F", x"0F", x"07", x"00", x"00", x"00", x"00", x"00", x"60", x"40", x"00", x"00", x"00", x"00", x"38", x"7C", x"9E", x"BE", x"FE", x"FE", x"7C", x"38", x"00", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"5C", x"7C", x"7C", x"38", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"30", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"56", x"56", x"7E", x"0D", x"00", x"00", x"00", x"3C", x"7E", x"7E", x"7E", x"FD", x"DB", x"FF", x"7E", x"3C", x"18", x"00", x"00", x"00", x"DB", x"FF", x"7E", x"3C", x"18", x"66", x"42", x"00", x"00", x"00", x"38", x"74", x"60", x"43", x"08", x"00", x"00", x"00", x"00", x"08", x"10", x"20", x"01", x"80", x"00", x"00", x"02", x"07", x"05", x"1F", x"07", x"01", x"00", x"03", x"05", x"00", x"00", x"1F", x"07", x"07", x"00", x"00", x"C0", x"E0", x"60", x"C0", x"80", x"F0", x"00", x"E0", x"30", x"10", x"10", x"30", x"F8", x"88", x"00", x"00", x"00", x"00", x"01", x"03", x"1F", x"00", x"07", x"07", x"07", x"07", x"06", x"0C", x"1F", x"00", x"F8", x"78", x"78", x"38", x"F8", x"F0", x"7C", x"00", x"00", x"80", x"80", x"C0", x"00", x"00", x"7C", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"FF", x"00", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"1C", x"0C", x"0E", x"07", x"03", x"01", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C3", x"FF", x"7E", x"00", x"FF", x"FF", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0E", x"0C", x"1C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"18", x"01", x"03", x"03", x"03", x"03", x"03", x"03", x"01", 
															x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"00", x"60", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"00", x"00", x"60", x"E0", x"C0", x"80", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7E", x"FE", x"C2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C3", x"81", x"00", x"00", x"00", x"00", x"81", x"C3", x"00", x"00", x"00", x"00", x"18", x"3C", x"7E", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"00", x"01", x"07", x"1F", x"7F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"00", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"39", x"39", x"1F", x"1F", x"0F", x"0F", x"04", x"00", x"46", x"46", x"20", x"20", x"10", x"10", x"0B", x"0C", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"00", x"B8", x"98", x"98", x"8C", x"8C", x"8C", x"00", x"00", x"00", x"60", x"20", x"10", x"10", x"10", x"C6", x"C6", x"C6", x"CE", x"D8", x"00", x"00", x"00", x"08", x"08", x"08", x"00", x"20", x"C0", x"00", x"00", x"00", x"F0", x"FE", x"FE", x"FE", x"FE", x"FC", x"CC", x"00", x"00", x"00", x"01", x"01", x"01", x"02", x"32", x"CC", x"F8", x"F8", x"F8", x"F0", x"F0", x"00", x"00", x"32", x"04", x"04", x"04", x"08", x"08", x"F8", x"00", 
															x"00", x"00", x"3E", x"30", x"30", x"30", x"30", x"30", x"00", x"00", x"01", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"07", x"0D", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"02", x"08", x"04", x"02", x"01", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"3E", x"1B", x"0E", x"04", x"00", x"00", x"00", x"00", x"40", x"24", x"11", x"0A", x"04", x"00", x"00", x"00", x"02", x"07", x"0D", x"07", x"13", x"21", x"40", x"C0", x"00", x"00", x"02", x"08", x"04", x"02", x"01", x"00", x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"1B", x"0E", x"04", x"08", x"10", x"A0", x"C0", x"40", x"24", x"11", x"0A", x"04", x"00", x"00", x"00", 
															x"00", x"80", x"C0", x"F0", x"F8", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"80", x"E0", x"F0", x"FC", x"FE", x"00", x"00", x"00", x"C0", x"E0", x"F8", x"FC", x"FF", x"00", x"00", x"00", x"00", x"80", x"C0", x"F0", x"F8", x"FF", x"FF", x"FF", x"FF", x"3F", x"07", x"00", x"00", x"FF", x"FF", x"FF", x"1F", x"03", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"1F", x"03", x"00", x"00", x"00", x"FE", x"7F", x"0F", x"01", x"00", x"00", x"00", x"00", x"80", x"E0", x"F0", x"F8", x"FC", x"7C", x"00", x"00", x"00", x"00", x"C0", x"E0", x"30", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"E0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F0", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"E0", x"00", x"00", x"FE", x"FF", x"FF", x"FE", x"F0", x"00", x"00", x"00", x"00", x"FE", x"FE", x"E0", x"00", x"00", x"00", x"00", 
															x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"3F", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"03", x"1F", x"FF", x"FF", x"03", x"1F", x"FF", x"FF", x"FF", x"FF", x"FC", x"F8", x"00", x"01", x"0F", x"7F", x"FE", x"F8", x"F0", x"C0", x"00", x"7C", x"FC", x"F8", x"F0", x"E0", x"80", x"00", x"00", x"00", x"30", x"E0", x"C0", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"F8", x"F0", x"C0", x"80", x"FF", x"FE", x"FC", x"F0", x"E0", x"80", x"00", x"00", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0E", x"1C", x"38", x"70", x"E0", x"C0", x"03", x"17", x"3E", x"7C", x"38", x"70", x"E0", x"C0", x"01", x"03", x"06", x"0C", x"18", x"30", x"60", x"C0", x"01", x"03", x"06", x"0C", x"18", x"30", x"60", x"C0", 
															x"00", x"01", x"03", x"05", x"07", x"1E", x"07", x"06", x"00", x"00", x"00", x"00", x"00", x"1F", x"07", x"01", x"00", x"00", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"E0", x"70", x"70", x"70", x"F0", x"F0", x"F0", x"2F", x"2F", x"2F", x"3F", x"1F", x"17", x"00", x"00", x"20", x"20", x"20", x"30", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"F8", x"F0", x"00", x"F8", x"FC", x"FE", x"F0", x"78", x"38", x"F0", x"00", x"00", x"00", x"01", x"03", x"02", x"03", x"02", x"07", x"00", x"03", x"06", x"24", x"24", x"35", x"3E", x"3F", x"00", x"00", x"40", x"E0", x"A0", x"E0", x"20", x"F0", x"00", x"E0", x"B0", x"12", x"12", x"D6", x"3E", x"FE", x"03", x"03", x"07", x"07", x"0F", x"07", x"00", x"00", x"1C", x"0C", x"0B", x"0F", x"06", x"06", x"00", x"00", x"E0", x"E0", x"F0", x"F0", x"E0", x"E0", x"F8", x"00", x"1C", x"18", x"08", x"08", x"10", x"60", x"F8", x"00", 
															x"00", x"00", x"01", x"03", x"03", x"01", x"00", x"00", x"00", x"03", x"06", x"04", x"04", x"06", x"07", x"0F", x"00", x"00", x"A0", x"F0", x"50", x"FC", x"F0", x"F0", x"00", x"E0", x"50", x"00", x"00", x"7C", x"F0", x"C8", x"00", x"01", x"01", x"01", x"01", x"03", x"1F", x"00", x"1F", x"3E", x"3E", x"26", x"06", x"04", x"1F", x"00", x"F8", x"F8", x"F8", x"F8", x"F8", x"F0", x"7C", x"00", x"04", x"04", x"06", x"02", x"00", x"00", x"7C", x"00", x"00", x"00", x"01", x"03", x"02", x"03", x"01", x"03", x"00", x"03", x"06", x"04", x"04", x"04", x"07", x"0F", x"00", x"00", x"40", x"E0", x"A0", x"E0", x"C0", x"E0", x"00", x"E0", x"B0", x"10", x"10", x"90", x"F0", x"F8", x"03", x"07", x"07", x"07", x"07", x"07", x"1F", x"00", x"0C", x"08", x"18", x"18", x"00", x"04", x"1F", x"00", x"E0", x"F0", x"F0", x"F0", x"F0", x"E0", x"78", x"00", x"18", x"08", x"0C", x"0C", x"00", x"20", x"78", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", x"00", x"01", x"0F", x"00", x"00", x"00", x"01", x"0F", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"38", x"E0", x"00", x"00", x"00", x"38", x"E0", x"00", x"00", x"00", x"00", x"80", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"0F", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"00", x"07", x"01", x"00", x"00", x"00", x"38", x"E0", x"00", x"00", x"00", x"00", x"80", x"F0", x"00", x"00", x"00", x"00", x"C0", x"70", x"00", x"03", x"0E", x"00", x"00", x"03", x"0E", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"00", x"07", x"38", x"E0", x"00", x"00", x"38", x"E0", x"00", x"00", x"00", x"00", x"00", x"F0", x"00", x"00", x"00", x"F0", 
															x"00", x"0F", x"00", x"00", x"0F", x"00", x"00", x"0F", x"00", x"00", x"07", x"00", x"00", x"07", x"00", x"00", x"F8", x"80", x"00", x"F8", x"80", x"00", x"F8", x"80", x"00", x"00", x"F0", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"0F", x"00", x"00", x"0F", x"00", x"00", x"07", x"00", x"00", x"07", x"00", x"00", x"07", x"00", x"00", x"F8", x"80", x"00", x"F8", x"80", x"00", x"F8", x"F0", x"00", x"00", x"F0", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"0F", x"00", x"00", x"0F", x"00", x"00", x"00", x"00", x"00", x"07", x"00", x"00", x"07", x"00", x"00", x"00", x"F8", x"00", x"F8", x"80", x"00", x"00", x"00", x"00", x"00", x"F0", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"6C", x"6C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"38", x"7C", x"FE", x"FE", x"FE", x"FE", x"7C", x"38", x"10", x"34", x"32", x"32", x"32", x"32", x"34", x"10", x"00", x"02", x"06", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"02", x"0E", x"08", x"08", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"02", x"0E", x"02", x"02", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"14", x"14", x"14", x"1E", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"08", x"0E", x"02", x"02", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"08", x"0E", x"0A", x"0A", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"0A", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"0E", x"0A", x"0E", x"0A", x"0A", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0E", x"0A", x"0E", x"02", x"02", x"0E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2E", x"6A", x"2A", x"2A", x"2A", x"2E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"3E", x"7F", x"7F", x"7F", x"7F", x"3E", x"1C", x"14", x"24", x"66", x"66", x"66", x"66", x"24", x"14", x"00", x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00", x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00", x"38", x"4C", x"18", x"30", x"60", x"7C", x"00", x"00", x"38", x"4C", x"18", x"30", x"60", x"7C", x"00", x"00", x"26", x"69", x"29", x"29", x"29", x"26", x"00", x"00", x"26", x"69", x"29", x"29", x"29", x"26", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"00", 
															x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"38", x"4C", x"C6", x"C6", x"C6", x"64", x"38", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"18", x"38", x"18", x"18", x"18", x"18", x"7E", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"7C", x"C6", x"0E", x"3C", x"78", x"E0", x"FE", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"7E", x"0C", x"18", x"3C", x"06", x"C6", x"7C", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"1C", x"3C", x"6C", x"CC", x"FE", x"0C", x"0C", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"FC", x"C0", x"FC", x"06", x"06", x"C6", x"7C", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"3C", x"60", x"C0", x"FC", x"C6", x"C6", x"7C", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", x"FE", x"C6", x"0C", x"18", x"30", x"30", x"30", x"00", 
															x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"7C", x"C6", x"C6", x"7C", x"C6", x"C6", x"7C", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"7C", x"C6", x"C6", x"7E", x"06", x"0C", x"78", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"38", x"6C", x"C6", x"C6", x"FE", x"C6", x"C6", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"FC", x"C6", x"C6", x"FC", x"C6", x"C6", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"1C", x"3C", x"1C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"60", x"70", x"78", x"70", x"60", x"40", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"FE", x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"8F", x"8F", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"7E", x"00", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", x"C6", x"E6", x"F6", x"FE", x"DE", x"CE", x"C6", x"00", 
															x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"7C", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"FC", x"C6", x"C6", x"C6", x"FC", x"C0", x"C0", x"00", x"8F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"FC", x"C6", x"C6", x"CE", x"F8", x"DC", x"CE", x"00", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"78", x"CC", x"C0", x"7C", x"06", x"C6", x"7C", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"7E", x"18", x"18", x"18", x"18", x"18", x"18", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"C6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7C", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"81", x"01", x"01", x"01", x"01", x"01", x"01", x"01", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"3E", x"60", x"C0", x"CE", x"C6", x"66", x"3E", x"00", x"38", x"7C", x"9E", x"BE", x"FE", x"FE", x"7C", x"38", x"38", x"7C", x"FE", x"FE", x"FE", x"FE", x"7C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"78", x"E0", x"C0", x"80", x"00", x"00", x"00", x"3C", x"78", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"60", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"60", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"70", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"70", 
															x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"80", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"80", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"3F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"60", x"40", x"40", x"40", x"40", x"40", x"4F", x"FC", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"06", x"02", x"02", x"02", x"02", x"02", x"F2", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"4F", x"49", x"48", x"48", x"48", x"49", x"49", x"4F", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"F2", x"92", x"92", x"12", x"12", x"12", x"92", x"F2", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"4F", x"40", x"40", x"40", x"40", x"40", x"60", x"3F", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"F2", x"02", x"02", x"02", x"02", x"02", x"06", x"FC", 
															x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FC", x"00", x"00", x"00", x"00", x"00", x"01", x"07", x"0C", x"FF", x"FF", x"FF", x"FC", x"F0", x"C0", x"00", x"00", x"00", x"01", x"07", x"1C", x"70", x"C0", x"00", x"00", x"FF", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"3F", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"0F", x"01", x"00", x"00", x"00", x"00", x"00", x"F8", x"0F", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"3F", x"0F", x"03", x"00", x"00", x"00", x"00", x"E0", x"38", x"0E", x"03", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"00", x"00", x"00", x"00", x"00", x"80", x"E0", x"30", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F8", x"00", x"00", x"00", x"01", x"03", x"06", x"0C", x"18", x"F8", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"38", x"60", x"C0", x"80", x"00", x"00", x"00", x"00", x"1F", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"1C", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"3F", x"1F", x"00", x"00", x"00", x"80", x"C0", x"60", x"30", x"18", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"F0", x"F0", x"E0", x"C0", x"C0", x"80", x"00", x"00", x"10", x"30", x"60", x"40", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"3F", x"7F", x"FF", x"00", x"00", x"00", x"03", x"0E", x"38", x"60", x"C0", 
															x"00", x"00", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"00", x"00", x"E0", x"B0", x"18", x"0C", x"06", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0F", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"F0", x"E0", x"C0", x"80", x"00", x"00", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"01", x"03", x"06", x"0C", x"18", x"30", x"60", x"C0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"FC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E0", x"3C", x"07", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"FC", x"FE", x"FF", x"00", x"00", x"00", x"C0", x"70", x"1C", x"06", x"03", x"0F", x"0F", x"07", x"03", x"03", x"01", x"00", x"00", x"08", x"0C", x"06", x"02", x"03", x"01", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"90", x"90", x"90", x"90", x"90", x"90", x"90", x"90", x"FE", x"FE", x"FC", x"FC", x"F8", x"F8", x"F0", x"F0", x"02", x"06", x"04", x"0C", x"08", x"18", x"10", x"10", x"01", x"01", x"03", x"07", x"07", x"0F", x"0F", x"1F", x"01", x"01", x"03", x"06", x"04", x"0C", x"08", x"18", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F0", x"F8", x"FC", x"FE", x"FF", x"80", x"C0", x"60", x"30", x"18", x"0C", x"06", x"03", x"00", x"00", x"00", x"00", x"18", x"3C", x"7E", x"FF", x"00", x"00", x"00", x"00", x"18", x"3C", x"66", x"C3", 
															x"80", x"80", x"C0", x"E0", x"E0", x"F0", x"F8", x"F8", x"80", x"80", x"C0", x"60", x"20", x"30", x"18", x"08", x"7F", x"7F", x"3F", x"3F", x"1F", x"1F", x"0F", x"0F", x"40", x"60", x"20", x"30", x"10", x"18", x"08", x"0C", x"F0", x"E0", x"E0", x"E0", x"C0", x"C0", x"C0", x"C0", x"30", x"20", x"20", x"60", x"40", x"40", x"40", x"C0", x"1F", x"3F", x"3F", x"7F", x"7F", x"7F", x"FF", x"FF", x"10", x"30", x"20", x"60", x"40", x"40", x"C0", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"00", x"00", x"00", x"07", x"1F", x"3F", x"7F", x"7F", x"00", x"00", x"00", x"00", x"00", x"C0", x"F0", x"F8", x"00", x"00", x"00", x"E0", x"F8", x"FC", x"FE", x"FE", 
															x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"FC", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"0C", x"04", x"06", x"02", x"02", x"03", x"01", x"01", x"07", x"07", x"07", x"03", x"03", x"03", x"03", x"01", x"04", x"04", x"06", x"02", x"02", x"02", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"1F", x"36", x"25", x"35", x"35", x"35", x"36", x"1F", x"FF", x"F6", x"E5", x"F5", x"F5", x"F5", x"F6", x"FF", x"F8", x"EC", x"54", x"54", x"54", x"54", x"EC", x"F8", x"FF", x"EF", x"57", x"57", x"57", x"57", x"EF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FC", x"F0", x"E0", x"C0", x"80", x"00", x"01", x"07", x"1C", x"30", x"60", x"C0", x"80", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"3F", x"0F", x"07", x"03", x"01", x"00", x"00", x"E0", x"38", x"0C", x"06", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"C0", x"E0", x"80", x"80", x"80", x"C0", x"40", x"40", x"40", x"60", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", 
															x"00", x"EE", x"AA", x"AA", x"AA", x"AA", x"EE", x"00", x"00", x"EE", x"AA", x"AA", x"AA", x"AA", x"EE", x"00", x"FF", x"FE", x"FC", x"F8", x"F0", x"E0", x"C0", x"80", x"03", x"06", x"0C", x"18", x"30", x"60", x"C0", x"80", x"00", x"00", x"07", x"08", x"10", x"10", x"20", x"20", x"00", x"00", x"07", x"0F", x"1F", x"1F", x"3F", x"3F", x"00", x"00", x"E0", x"10", x"08", x"08", x"04", x"04", x"00", x"00", x"E0", x"F0", x"F8", x"F8", x"FC", x"FC", x"FF", x"FF", x"7F", x"7F", x"3F", x"3F", x"1F", x"1F", x"80", x"C0", x"40", x"60", x"20", x"30", x"10", x"18", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"80", x"80", x"80", x"C0", x"C0", x"C0", x"E0", x"E0", x"80", x"80", x"80", x"C0", x"40", x"40", x"60", x"20", x"FF", x"FF", x"FF", x"7F", x"7F", x"7F", x"3F", x"3F", x"80", x"80", x"C0", x"40", x"40", x"60", x"20", x"20", 
															x"20", x"20", x"10", x"10", x"08", x"07", x"00", x"00", x"3F", x"3F", x"1F", x"1F", x"0F", x"07", x"00", x"00", x"04", x"04", x"08", x"08", x"10", x"E0", x"00", x"00", x"FC", x"FC", x"F8", x"F8", x"F0", x"E0", x"00", x"00", x"00", x"0E", x"08", x"0E", x"02", x"02", x"0E", x"00", x"00", x"0E", x"08", x"0E", x"02", x"02", x"0E", x"00", x"00", x"2E", x"6A", x"2A", x"2A", x"2A", x"2E", x"00", x"00", x"2E", x"6A", x"2A", x"2A", x"2A", x"2E", x"00", x"0F", x"0F", x"0F", x"0F", x"07", x"07", x"07", x"07", x"08", x"08", x"08", x"0C", x"04", x"04", x"04", x"04", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"E0", x"F0", x"F0", x"F0", x"F8", x"F8", x"F8", x"FC", x"20", x"30", x"10", x"10", x"18", x"08", x"08", x"0C", x"3F", x"1F", x"1F", x"1F", x"0F", x"0F", x"0F", x"07", x"30", x"10", x"10", x"18", x"08", x"08", x"0C", x"04", 
															x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"01", x"C0", x"60", x"30", x"18", x"0C", x"06", x"03", x"01", x"01", x"03", x"07", x"0F", x"1F", x"3F", x"7F", x"FF", x"01", x"03", x"07", x"0D", x"19", x"31", x"61", x"C1", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"FC", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"04", x"04", x"06", x"02", x"02", x"03", x"01", x"01", x"07", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"06", x"02", x"03", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"7C", x"01", x"01", x"01", x"01", x"83", x"82", x"C6", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", 
															x"00", x"00", x"00", x"00", x"03", x"0F", x"1F", x"3F", x"0F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"C0", x"F0", x"F8", x"FC", x"F0", x"FC", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"07", x"07", x"07", x"07", x"07", x"03", x"3F", x"76", x"65", x"75", x"75", x"75", x"76", x"3F", x"FF", x"F6", x"E5", x"F5", x"F5", x"F5", x"F6", x"FF", x"FC", x"EE", x"56", x"56", x"56", x"56", x"EE", x"FC", x"FF", x"EF", x"57", x"57", x"57", x"57", x"EF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"01", x"01", x"00", x"00", x"00", x"00", 
															x"3F", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", x"3F", x"0F", x"FC", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"60", x"60", x"60", x"60", x"60", x"00", x"07", x"07", x"07", x"0F", x"0F", x"0F", x"1F", x"1F", x"04", x"04", x"04", x"0C", x"08", x"08", x"18", x"10", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"06", x"1F", x"3F", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"10", x"30", x"20", x"60", x"C0", x"80", x"00", x"00", x"0F", x"3F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"0C", x"38", x"E0", x"80", x"80", x"80", x"80", x"80", 
															x"00", x"00", x"00", x"03", x"07", x"06", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"06", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"03", x"03", x"C0", x"60", x"30", x"18", x"0C", x"06", x"02", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"1C", x"1E", x"1B", x"19", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D8", x"D8", x"C0", x"DA", x"DB", x"DB", x"DB", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"1E", x"CC", x"6D", x"6D", x"6D", x"6C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E5", x"B6", x"F6", x"86", x"E6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"8F", x"DB", x"DB", x"DB", x"CF", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"6C", x"6C", x"6C", x"38", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"01", x"03", x"07", x"07", x"07", x"07", x"07", x"07", x"01", x"03", x"06", x"04", x"04", x"04", x"04", x"04", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"F8", x"FF", x"FF", x"FF", x"FF", x"80", x"C0", x"60", x"38", x"0F", x"00", x"00", x"00", x"03", x"07", x"0F", x"3F", x"FF", x"FF", x"FF", x"FF", x"02", x"06", x"0C", x"38", x"E0", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", 
															x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"FF", x"FF", x"FE", x"FE", x"FC", x"FC", x"F8", x"F8", x"01", x"03", x"02", x"06", x"04", x"0C", x"08", x"18", x"1F", x"0F", x"03", x"00", x"00", x"00", x"00", x"00", x"7F", x"7F", x"3F", x"1F", x"07", x"00", x"00", x"00", x"F8", x"F0", x"C0", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FC", x"F8", x"E0", x"00", x"00", x"00", x"0F", x"0F", x"07", x"07", x"03", x"03", x"01", x"01", x"08", x"0C", x"04", x"06", x"02", x"03", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"3F", x"7F", x"5B", x"55", x"55", x"55", x"5B", x"7F", x"3F", x"7F", x"5B", x"55", x"55", x"55", x"5B", x"7F", x"FC", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", 
															x"3F", x"7F", x"63", x"77", x"77", x"57", x"67", x"7F", x"3F", x"7F", x"63", x"77", x"77", x"57", x"67", x"7F", x"3F", x"7F", x"67", x"5B", x"5B", x"57", x"63", x"7F", x"3F", x"7F", x"67", x"5B", x"5B", x"57", x"63", x"7F", x"3F", x"7F", x"5B", x"57", x"4F", x"57", x"5B", x"7F", x"3F", x"7F", x"5B", x"57", x"4F", x"57", x"5B", x"7F", x"3F", x"7F", x"67", x"5B", x"5B", x"43", x"5B", x"7F", x"3F", x"7F", x"67", x"5B", x"5B", x"43", x"5B", x"7F", x"7F", x"7F", x"7E", x"7C", x"7C", x"7F", x"7E", x"7F", x"7F", x"7F", x"7E", x"7C", x"7C", x"7F", x"7E", x"7F", x"FE", x"7E", x"3E", x"1E", x"9E", x"7E", x"3E", x"FE", x"FE", x"7E", x"3E", x"1E", x"9E", x"7E", x"3E", x"FE", x"0F", x"07", x"03", x"03", x"01", x"01", x"01", x"01", x"0C", x"06", x"02", x"03", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"03", x"07", x"07", x"0F", x"01", x"01", x"01", x"03", x"02", x"06", x"04", x"0C", 
															x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"3F", x"FE", x"DA", x"AA", x"AA", x"AA", x"DA", x"FE", x"FC", x"FE", x"DA", x"AA", x"AA", x"AA", x"DA", x"FE", x"FC", x"FE", x"E6", x"EA", x"EE", x"EE", x"C6", x"FE", x"FC", x"FE", x"E6", x"EA", x"EE", x"EE", x"C6", x"FE", x"FC", x"FE", x"C6", x"EA", x"DA", x"DA", x"E6", x"FE", x"FC", x"FE", x"C6", x"EA", x"DA", x"DA", x"E6", x"FE", x"FC", x"FE", x"DA", x"EA", x"F2", x"EA", x"DA", x"FE", x"FC", x"FE", x"DA", x"EA", x"F2", x"EA", x"DA", x"FE", x"FC", x"FE", x"DA", x"C2", x"DA", x"DA", x"E6", x"FE", x"FC", x"FE", x"DA", x"C2", x"DA", x"DA", x"E6", x"FE", x"FC", x"0F", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"FF", x"08", x"18", x"10", x"30", x"20", x"60", x"40", x"C0", x"00", x"FF", x"C5", x"DD", x"C6", x"DD", x"C5", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"00", x"FF", x"51", x"5B", x"DB", x"5B", x"5B", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"07", x"05", x"05", x"04", x"04", x"04", x"04", x"02", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"02", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"03", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"00", x"80", x"80", x"80", x"C0", x"40", x"00", x"00", x"00", x"80", x"80", x"80", x"C0", x"C0", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
															x"02", x"06", x"04", x"04", x"0C", x"08", x"08", x"18", x"03", x"07", x"07", x"07", x"0F", x"0F", x"0F", x"1F", x"40", x"E0", x"A0", x"A0", x"20", x"20", x"20", x"20", x"40", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"40", x"60", x"20", x"20", x"30", x"10", x"10", x"18", x"C0", x"E0", x"E0", x"E0", x"F0", x"F0", x"F0", x"F8", x"04", x"04", x"04", x"04", x"06", x"02", x"03", x"01", x"07", x"07", x"07", x"07", x"07", x"03", x"03", x"01", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"10", x"10", x"30", x"20", x"20", x"60", x"40", x"41", x"1F", x"1F", x"3F", x"3F", x"3F", x"7F", x"7F", x"7F", x"FF", x"FF", x"FF", x"FF", x"E6", x"E3", x"E0", x"E0", x"00", x"00", x"00", x"00", x"06", x"03", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"03", x"83", x"C3", x"73", x"00", x"00", x"00", x"00", x"00", x"80", x"C0", x"70", 
															x"03", x"03", x"03", x"03", x"03", x"01", x"01", x"00", x"03", x"03", x"03", x"03", x"03", x"01", x"01", x"00", x"08", x"08", x"0C", x"04", x"04", x"06", x"02", x"82", x"F8", x"F8", x"FC", x"FC", x"FC", x"FE", x"FE", x"FE", x"C3", x"71", x"1B", x"0E", x"00", x"00", x"00", x"00", x"FF", x"7F", x"1F", x"0E", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"20", x"60", x"40", x"C0", x"80", x"E0", x"E0", x"E0", x"E0", x"E0", x"C0", x"C0", x"80", x"C3", x"8E", x"D8", x"70", x"00", x"00", x"00", x"00", x"FF", x"FE", x"F8", x"70", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"80", x"80", x"00", x"E0", x"E0", x"E0", x"E0", x"E6", x"E3", x"E0", x"E0", x"00", x"00", x"03", x"0E", x"06", x"03", x"00", x"00", x"00", x"03", x"03", x"03", x"03", x"83", x"C3", x"73", x"38", x"E0", x"80", x"00", x"00", x"80", x"C0", x"70", 
															x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"00", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"E0", x"70", x"3C", x"1E", x"07", x"03", x"01", x"00", x"E0", x"70", x"3C", x"1E", x"07", x"03", x"01", x"00", x"07", x"0E", x"3C", x"78", x"E0", x"C0", x"80", x"00", x"07", x"0E", x"3C", x"78", x"E0", x"C0", x"80", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"00", x"00", x"00", x"00", x"01", x"01", x"03", x"03", x"3C", x"1E", x"07", x"03", x"01", x"00", x"00", x"00", x"3C", x"1E", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0E", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0E", x"3F", x"60", x"C0", x"80", x"80", x"80", x"80", x"C0", x"3F", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"61", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", x"7F", x"3F", x"00", x"00", x"00", x"00", x"00", x"00", 
															x"FF", x"FD", x"FD", x"FF", x"FF", x"FD", x"FD", x"FF", x"07", x"05", x"05", x"07", x"07", x"05", x"05", x"07", x"FF", x"99", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"99", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"BF", x"BF", x"FF", x"FF", x"BF", x"BF", x"FF", x"E0", x"A0", x"A0", x"E0", x"E0", x"A0", x"A0", x"E0", x"00", x"00", x"00", x"00", x"00", x"FF", x"99", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"99", x"FF", x"F0", x"F0", x"E0", x"E0", x"C0", x"C0", x"80", x"80", x"10", x"30", x"20", x"60", x"40", x"C0", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"0E", x"1F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"38", x"38", x"3C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"0F", x"0F", x"07", x"03", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"38", x"38", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0E", x"0C", x"1F", x"1F", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"F0", x"38", x"98", x"9C", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1E", x"0C", x"0C", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"18", x"18", x"F0", x"E0", x"00", x"00", x"00", x"80", x"80", x"C0", x"C0", x"E0", x"E0", x"F0", x"F0", x"80", x"80", x"C0", x"40", x"60", x"20", x"30", x"10", x"3E", x"63", x"C0", x"80", x"80", x"80", x"80", x"C0", x"3E", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"60", x"38", x"0F", x"01", x"00", x"00", x"00", x"00", x"7F", x"3F", x"0F", x"01", x"00", x"00", x"00", x"00", 
															x"01", x"01", x"03", x"03", x"07", x"07", x"0F", x"0F", x"01", x"01", x"03", x"02", x"06", x"04", x"0C", x"08", x"F8", x"F8", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"18", x"08", x"0C", x"04", x"06", x"02", x"03", x"01", x"F8", x"F8", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"18", x"08", x"0C", x"04", x"06", x"02", x"03", x"FF", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"FF", x"FF", x"18", x"10", x"30", x"20", x"60", x"40", x"C0", x"FF", x"1F", x"1F", x"3F", x"3F", x"7F", x"7F", x"FF", x"FF", x"18", x"10", x"30", x"20", x"60", x"40", x"C0", x"80", x"00", x"7F", x"3F", x"1F", x"07", x"03", x"01", x"FF", x"FF", x"FE", x"FC", x"F8", x"E0", x"C0", x"80", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"66", x"66", x"66", x"3C", x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1D", x"0C", x"0F", x"07", x"03", x"00", x"00", x"00", 
															x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"18", x"38", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1F", x"0C", x"0E", x"07", x"03", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"9C", x"98", x"38", x"F0", x"E0", x"00", x"00", x"00", x"00", x"00", x"01", x"03", x"07", x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"07", x"0F", x"0E", x"1D", x"1D", x"92", x"54", x"38", x"FE", x"38", x"54", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"0F", x"38", x"00", x"00", x"00", x"00", x"00", x"01", x"0F", x"3F", x"60", x"C0", x"80", x"80", x"80", x"80", x"C0", x"63", x"7F", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"7F", 
															x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"F0", x"1C", x"00", x"00", x"00", x"00", x"00", x"80", x"F0", x"FC", x"06", x"03", x"01", x"01", x"01", x"01", x"03", x"C6", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FC", x"06", x"03", x"01", x"01", x"01", x"01", x"03", x"FC", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"86", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"7C", x"C6", x"03", x"01", x"01", x"01", x"01", x"03", x"7C", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"06", x"1C", x"F0", x"80", x"00", x"00", x"00", x"00", x"FE", x"FC", x"F0", x"80", x"00", x"00", x"00", x"00");

END PACKAGE;