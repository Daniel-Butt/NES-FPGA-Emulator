library ieee;
use ieee.std_logic_1164.all;


PACKAGE opcodes IS

	CONSTANT BRK_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"00";
	CONSTANT ORA_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"01";
	CONSTANT ORA_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"05";
	CONSTANT ASL_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"06";
	CONSTANT PHP_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"08";
	CONSTANT ORA_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"09";
	CONSTANT ASL_A : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0a";
	CONSTANT ORA_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0d";
	CONSTANT ASL_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"0e";
	CONSTANT BPL_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"10";
	CONSTANT ORA_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"11";
	CONSTANT ORA_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"15";
	CONSTANT ASL_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"16";
	CONSTANT CLC_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"18";
	CONSTANT ORA_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"19";
	CONSTANT ORA_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1d";
	CONSTANT ASL_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"1e";
	CONSTANT JSR_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"20";
	CONSTANT AND_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"21";
	CONSTANT BIT_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"24";
	CONSTANT AND_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"25";
	CONSTANT ROL_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"26";
	CONSTANT PLP_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"28";
	CONSTANT AND_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"29";
	CONSTANT ROL_A : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"2a";
	CONSTANT BIT_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"2c";
	CONSTANT AND_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"2d";
	CONSTANT ROL_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"2e";
	CONSTANT BMI_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"30";
	CONSTANT AND_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"31";
	CONSTANT AND_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"35";
	CONSTANT ROL_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"36";
	CONSTANT SEC_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"38";
	CONSTANT AND_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"39";
	CONSTANT AND_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"3d";
	CONSTANT ROL_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"3e";
	CONSTANT RTI_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"40";
	CONSTANT EOR_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"41";
	CONSTANT EOR_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"45";
	CONSTANT LSR_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"46";
	CONSTANT PHA_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"48";
	CONSTANT EOR_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"49";
	CONSTANT LSR_A : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"4a";
	CONSTANT JMP_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"4c";
	CONSTANT EOR_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"4d";
	CONSTANT LSR_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"4e";
	CONSTANT BVC_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"50";
	CONSTANT EOR_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"51";
	CONSTANT EOR_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"55";
	CONSTANT LSR_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"56";
	CONSTANT CLI_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"58";
	CONSTANT EOR_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"59";
	CONSTANT EOR_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"5d";
	CONSTANT LSR_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"5e";
	CONSTANT RTS_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"60";
	CONSTANT ADC_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"61";
	CONSTANT ADC_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"65";
	CONSTANT ROR_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"66";
	CONSTANT PLA_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"68";
	CONSTANT ADC_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"69";
	CONSTANT ROR_A : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"6a";
	CONSTANT JMP_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"6c";
	CONSTANT ADC_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"6d";
	CONSTANT ROR_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"6e";
	CONSTANT BVS_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"70";
	CONSTANT ADC_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"71";
	CONSTANT ADC_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"75";
	CONSTANT ROR_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"76";
	CONSTANT SEI_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"78";
	CONSTANT ADC_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"79";
	CONSTANT ADC_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"7d";
	CONSTANT ROR_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"7e";
	CONSTANT STA_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"81";
	CONSTANT STY_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"84";
	CONSTANT STA_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"85";
	CONSTANT STX_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"86";
	CONSTANT DEY_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"88";
	CONSTANT TXA_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"8a";
	CONSTANT STY_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"8c";
	CONSTANT STA_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"8d";
	CONSTANT STX_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"8e";
	CONSTANT BCC_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"90";
	CONSTANT STA_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"91";
	CONSTANT STY_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"94";
	CONSTANT STA_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"95";
	CONSTANT STX_ZPG_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"96";
	CONSTANT TYA_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"98";
	CONSTANT STA_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"99";
	CONSTANT TXS_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"9a";
	CONSTANT STA_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"9d";
	CONSTANT LDY_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a0";
	CONSTANT LDA_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a1";
	CONSTANT LDX_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a2";
	CONSTANT LDY_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a4";
	CONSTANT LDA_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a5";
	CONSTANT LDX_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a6";
	CONSTANT TAY_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a8";
	CONSTANT LDA_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"a9";
	CONSTANT TAX_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"aa";
	CONSTANT LDY_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ac";
	CONSTANT LDA_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ad";
	CONSTANT LDX_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ae";
	CONSTANT BCS_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b0";
	CONSTANT LDA_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b1";
	CONSTANT LDY_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b4";
	CONSTANT LDA_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b5";
	CONSTANT LDX_ZPG_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b6";
	CONSTANT CLV_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b8";
	CONSTANT LDA_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"b9";
	CONSTANT TSX_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ba";
	CONSTANT LDY_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"bc";
	CONSTANT LDA_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"bd";
	CONSTANT LDX_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"be";
	CONSTANT CPY_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c0";
	CONSTANT CMP_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c1";
	CONSTANT CPY_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c4";
	CONSTANT CMP_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c5";
	CONSTANT DEC_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c6";
	CONSTANT INY_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c8";
	CONSTANT CMP_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"c9";
	CONSTANT DEX_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ca";
	CONSTANT CPY_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"cc";
	CONSTANT CMP_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"cd";
	CONSTANT DEC_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ce";
	CONSTANT BNE_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"d0";
	CONSTANT CMP_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"d1";
	CONSTANT CMP_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"d5";
	CONSTANT DEC_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"d6";
	CONSTANT CLD_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"d8";
	CONSTANT CMP_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"d9";
	CONSTANT CMP_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"dd";
	CONSTANT DEC_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"de";
	CONSTANT CPX_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e0";
	CONSTANT SBC_X_IND : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e1";
	CONSTANT CPX_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e4";
	CONSTANT SBC_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e5";
	CONSTANT INC_ZPG : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e6";
	CONSTANT INX_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e8";
	CONSTANT SBC_IMM : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"e9";
	CONSTANT NOP_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ea";
	CONSTANT CPX_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ec";
	CONSTANT SBC_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ed";
	CONSTANT INC_ABS : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"ee";
	CONSTANT BEQ_REL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"f0";
	CONSTANT SBC_IND_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"f1";
	CONSTANT SBC_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"f5";
	CONSTANT INC_ZPG_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"f6";
	CONSTANT SED_IMPL : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"f8";
	CONSTANT SBC_ABS_Y : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"f9";
	CONSTANT SBC_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"fd";
	CONSTANT INC_ABS_X : STD_LOGIC_VECTOR(7 DOWNTO 0) :=x"fe";


END PACKAGE;